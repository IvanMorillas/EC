//: version "1.8.7"

module sumador_HA2(S, C, Cin, B, A);
//: interface  /sz:(172, 140) /bd:[ Li0>Cin(106/140) Li1>B(68/140) Li2>A(29/140) Ro0<C(82/140) Ro1<S(44/140) ]
input B;    //: /sn:0 {0}(364,208)(364,258){1}
//: {2}(366,260)(454,260)(454,256)(613,256){3}
//: {4}(364,262)(364,391){5}
//: {6}(366,393)(543,393){7}
//: {8}(364,395)(364,415)(543,415){9}
input A;    //: /sn:0 {0}(544,361)(325,361){1}
//: {2}(323,359)(323,253){3}
//: {4}(325,251)(613,251){5}
//: {6}(323,249)(323,209){7}
//: {8}(323,363)(323,379)(335,379)(335,388)(543,388){9}
input Cin;    //: /sn:0 /dp:3 {0}(398,210)(398,270){1}
//: {2}(400,272)(498,272)(498,267)(732,267){3}
//: {4}(398,274)(398,363){5}
//: {6}(400,365)(410,365)(410,366)(544,366){7}
//: {8}(398,367)(398,420)(543,420){9}
output C;    //: /sn:0 {0}(1031,318)(811,318)(811,317)(810,317){1}
output S;    //: /sn:0 /dp:1 {0}(753,265)(1025,265)(1025,251)(1035,251){1}
wire w16;    //: /sn:0 /dp:1 {0}(692,322)(654,322)(654,391)(564,391){1}
wire w8;    //: /sn:0 {0}(564,418)(779,418)(779,319)(789,319){1}
wire w11;    //: /sn:0 {0}(634,254)(722,254)(722,262)(732,262){1}
wire w15;    //: /sn:0 /dp:1 {0}(692,317)(626,317)(626,364)(565,364){1}
wire w5;    //: /sn:0 /dp:1 {0}(789,314)(735,314)(735,320)(713,320){1}
//: enddecls

  //: output g4 (S) @(1032,251) /sn:0 /w:[ 1 ]
  xor g8 (.I0(A), .I1(B), .Z(w11));   //: @(624,254) /sn:0 /delay:" 4" /w:[ 5 3 0 ]
  //: output g3 (C) @(1028,318) /sn:0 /w:[ 0 ]
  //: joint g16 (Cin) @(398, 365) /w:[ 6 5 -1 8 ]
  //: input g2 (Cin) @(398,208) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (B) @(364,206) /sn:0 /R:3 /w:[ 0 ]
  //: joint g18 (B) @(364, 393) /w:[ 6 5 -1 8 ]
  or g10 (.I0(w15), .I1(w16), .Z(w5));   //: @(703,320) /sn:0 /delay:" 3" /w:[ 0 0 1 ]
  and g6 (.I0(A), .I1(B), .Z(w16));   //: @(554,391) /sn:0 /delay:" 3" /w:[ 9 7 1 ]
  and g7 (.I0(B), .I1(Cin), .Z(w8));   //: @(554,418) /sn:0 /delay:" 3" /w:[ 9 9 0 ]
  xor g9 (.I0(w11), .I1(Cin), .Z(S));   //: @(743,265) /sn:0 /delay:" 4" /w:[ 1 3 0 ]
  //: joint g12 (A) @(323, 251) /w:[ 4 6 -1 3 ]
  and g5 (.I0(A), .I1(Cin), .Z(w15));   //: @(555,364) /sn:0 /delay:" 3" /w:[ 0 7 1 ]
  or g11 (.I0(w5), .I1(w8), .Z(C));   //: @(800,317) /sn:0 /delay:" 3" /w:[ 0 1 1 ]
  //: joint g14 (Cin) @(398, 272) /w:[ 2 1 -1 4 ]
  //: input g0 (A) @(323,207) /sn:0 /R:3 /w:[ 7 ]
  //: joint g15 (A) @(323, 361) /w:[ 1 2 -1 8 ]
  //: joint g13 (B) @(364, 260) /w:[ 2 1 -1 4 ]

endmodule

module CPA_2(Cin, A, B, S);
//: interface  /sz:(212, 165) /bd:[ Li0>A[3:0](36/165) Li1>B[3:0](77/165) Li2>Cin(121/165) Ro0<S[4:0](48/165) ]
input [3:0] B;    //: /sn:0 {0}(1126,100)(1025,100){1}
//: {2}(1024,100)(819,100){3}
//: {4}(818,100)(628,100){5}
//: {6}(627,100)(404,100){7}
//: {8}(403,100)(361,100){9}
input [3:0] A;    //: /sn:0 {0}(1075,60)(1065,60){1}
//: {2}(1064,60)(780,60){3}
//: {4}(779,60)(666,60){5}
//: {6}(665,60)(444,60){7}
//: {8}(443,60)(202,60){9}
input Cin;    //: /sn:0 /dp:1 {0}(971,185)(987,185)(987,206){1}
output [4:0] S;    //: /sn:0 /dp:1 {0}(1151,526)(1225,526)(1225,539)(1343,539){1}
wire w6;    //: /sn:0 {0}(629,209)(629,112)(628,112)(628,104){1}
wire w16;    //: /sn:0 {0}(1025,206)(1025,104){1}
wire w13;    //: /sn:0 {0}(834,380)(834,390)(717,390)(717,199)(591,199)(591,209){1}
wire w7;    //: /sn:0 {0}(668,209)(668,72)(666,72)(666,64){1}
wire w4;    //: /sn:0 {0}(429,387)(429,516)(1145,516){1}
wire w3;    //: /sn:0 {0}(391,387)(391,506)(1145,506){1}
wire w12;    //: /sn:0 /dp:1 {0}(781,206)(781,68)(780,68)(780,64){1}
wire w19;    //: /sn:0 {0}(1049,380)(1049,546)(1145,546){1}
wire w18;    //: /sn:0 {0}(1011,380)(1011,390)(926,390)(926,196)(858,196)(858,206){1}
wire w1;    //: /sn:0 {0}(405,213)(405,112)(404,112)(404,104){1}
wire w8;    //: /sn:0 {0}(615,383)(615,393)(515,393)(515,203)(367,203)(367,213){1}
wire w17;    //: /sn:0 {0}(1064,206)(1064,72)(1065,72)(1065,64){1}
wire w14;    //: /sn:0 {0}(796,380)(796,536)(1145,536){1}
wire w2;    //: /sn:0 {0}(444,213)(444,64){1}
wire w11;    //: /sn:0 {0}(820,206)(820,112)(819,112)(819,104){1}
wire w9;    //: /sn:0 {0}(653,383)(653,526)(1145,526){1}
//: enddecls

  tran g8(.Z(w17), .I(A[0]));   //: @(1065,58) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: input g4 (Cin) @(969,185) /sn:0 /w:[ 0 ]
  tran g16(.Z(w1), .I(B[3]));   //: @(404,98) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  sumador_HA2 g3 (.A(w17), .B(w16), .Cin(Cin), .S(w19), .C(w18));   //: @(953, 207) /sz:(140, 172) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  sumador_HA2 g2 (.A(w12), .B(w11), .Cin(w18), .S(w14), .C(w13));   //: @(752, 207) /sz:(140, 172) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  sumador_HA2 g1 (.A(w7), .B(w6), .Cin(w13), .S(w9), .C(w8));   //: @(557, 210) /sz:(140, 172) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  tran g10(.Z(w7), .I(A[2]));   //: @(666,58) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  concat g6 (.I0(w19), .I1(w14), .I2(w9), .I3(w4), .I4(w3), .Z(S));   //: @(1150,526) /sn:0 /w:[ 1 1 1 1 1 0 ] /dr:0
  tran g9(.Z(w12), .I(A[1]));   //: @(780,58) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: input g7 (A) @(200,60) /sn:0 /w:[ 9 ]
  //: input g12 (B) @(1128,100) /sn:0 /R:2 /w:[ 0 ]
  tran g14(.Z(w11), .I(B[1]));   //: @(819,98) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g11(.Z(w2), .I(A[3]));   //: @(444,58) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  //: output g5 (S) @(1340,539) /sn:0 /w:[ 1 ]
  tran g15(.Z(w6), .I(B[2]));   //: @(628,98) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  sumador_HA2 g0 (.A(w2), .B(w1), .Cin(w8), .S(w4), .C(w3));   //: @(333, 214) /sz:(140, 172) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  tran g13(.Z(w16), .I(B[0]));   //: @(1025,98) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1

endmodule

module main;    //: root_module
wire [3:0] w4;    //: /sn:0 {0}(294,322)(294,352)(487,352){1}
wire [4:0] w0;    //: /sn:0 {0}(701,323)(933,323)(933,236){1}
wire [3:0] w1;    //: /sn:0 /dp:1 {0}(487,311)(382,311)(382,298){1}
wire w2;    //: /sn:0 {0}(414,396)(487,396){1}
//: enddecls

  led g4 (.I(w0));   //: @(933,229) /sn:0 /w:[ 1 ] /type:3
  //: switch g3 (w2) @(397,396) /sn:0 /w:[ 0 ] /st:0
  //: dip g2 (w4) @(294,312) /sn:0 /w:[ 0 ] /st:0
  //: dip g1 (w1) @(382,288) /sn:0 /w:[ 1 ] /st:0
  CPA_2 g0 (.Cin(w2), .B(w4), .A(w1), .S(w0));   //: @(488, 275) /sz:(212, 165) /sn:0 /p:[ Li0>1 Li1>1 Li2>0 Ro0<0 ]

endmodule
