//: version "1.8.7"

module Sumador_HA(C, B, A, S);
//: interface  /sz:(183, 129) /bd:[ Li0>A(35/129) Li1>B(80/129) Ro0<S(62/129) Ro1<C(89/129) ]
input B;    //: /sn:0 {0}(354,174)(393,174)(393,173)(403,173){1}
//: {2}(407,173)(424,173)(424,159)(432,159){3}
//: {4}(405,175)(405,193)(429,193){5}
input A;    //: /sn:0 {0}(353,155)(380,155)(380,154)(390,154){1}
//: {2}(394,154)(432,154){3}
//: {4}(392,156)(392,188)(429,188){5}
output C;    //: /sn:0 {0}(515,191)(450,191){1}
output S;    //: /sn:0 {0}(515,157)(453,157){1}
//: enddecls

  //: output g4 (C) @(512,191) /sn:0 /w:[ 0 ]
  //: input g3 (B) @(352,174) /sn:0 /w:[ 0 ]
  //: input g2 (A) @(351,155) /sn:0 /w:[ 0 ]
  xor g1 (.I0(A), .I1(B), .Z(S));   //: @(443,157) /sn:0 /delay:" 4" /w:[ 3 3 1 ]
  //: joint g6 (A) @(392, 154) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(405, 173) /w:[ 2 -1 1 4 ]
  //: output g5 (S) @(512,157) /sn:0 /w:[ 0 ]
  and g0 (.I0(A), .I1(B), .Z(C));   //: @(440,191) /sn:0 /delay:" 3" /w:[ 5 5 1 ]

endmodule

module Sumador_FA(B, A, C, S, Cin);
//: interface  /sz:(90, 70) /bd:[ Li0>A(11/59) Li1>B(28/59) Li2>Cin(43/59) Ro0<S(15/59) Ro1<C(36/59) ]
input B;    //: /sn:0 {0}(67,222)(120,222)(120,219)(130,219){1}
input A;    //: /sn:0 /dp:1 {0}(69,193)(120,193)(120,194)(130,194){1}
input Cin;    //: /sn:0 {0}(71,286)(327,286)(327,261)(337,261){1}
output C;    //: /sn:0 {0}(574,310)(544,310)(544,309)(514,309){1}
output S;    //: /sn:0 /dp:1 {0}(443,251)(584,251)(584,253)(594,253){1}
wire w7;    //: /sn:0 {0}(443,266)(483,266)(483,306)(493,306){1}
wire w2;    //: /sn:0 {0}(213,209)(273,209)(273,236)(337,236){1}
wire w9;    //: /sn:0 /dp:1 {0}(493,311)(264,311)(264,224)(213,224){1}
//: enddecls

  //: input g4 (B) @(65,222) /sn:0 /w:[ 0 ]
  //: input g3 (A) @(67,193) /sn:0 /w:[ 0 ]
  or g2 (.I0(w7), .I1(w9), .Z(C));   //: @(504,309) /sn:0 /delay:" 3" /w:[ 1 0 1 ]
  Sumador_HA g1 (.B(Cin), .A(w2), .C(w7), .S(S));   //: @(338, 218) /sz:(104, 70) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: output g6 (C) @(571,310) /sn:0 /w:[ 0 ]
  //: output g7 (S) @(591,253) /sn:0 /w:[ 1 ]
  //: input g5 (Cin) @(69,286) /sn:0 /w:[ 0 ]
  Sumador_HA g0 (.B(B), .A(A), .C(w9), .S(w2));   //: @(131, 176) /sz:(81, 70) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]

endmodule

module main;    //: root_module
wire w3;    //: /sn:0 {0}(422,189)(355,189){1}
wire w0;    //: /sn:0 {0}(205,180)(263,180){1}
wire w1;    //: /sn:0 {0}(205,207)(253,207)(253,198)(263,198){1}
wire w2;    //: /sn:0 {0}(425,164)(355,164){1}
wire w5;    //: /sn:0 {0}(205,153)(253,153)(253,160)(263,160){1}
//: enddecls

  led g4 (.I(w2));   //: @(432,164) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: switch g3 (w1) @(188,207) /sn:0 /w:[ 0 ] /st:1
  //: switch g2 (w0) @(188,180) /sn:0 /w:[ 0 ] /st:1
  //: switch g1 (w5) @(188,153) /sn:0 /w:[ 0 ] /st:1
  led g5 (.I(w3));   //: @(429,189) /sn:0 /R:3 /w:[ 0 ] /type:0
  Sumador_FA g0 (.Cin(w1), .B(w0), .A(w5), .C(w3), .S(w2));   //: @(264, 147) /sz:(90, 70) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Ro0<1 Ro1<1 ]

endmodule
