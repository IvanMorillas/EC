//: version "1.8.7"

module Sumador_HA(C, B, A, S);
//: interface  /sz:(183, 129) /bd:[ Li0>A(35/129) Li1>B(80/129) Ro0<S(62/129) Ro1<C(89/129) ]
input B;    //: /sn:0 {0}(354,174)(393,174)(393,173)(403,173){1}
//: {2}(407,173)(424,173)(424,159)(432,159){3}
//: {4}(405,175)(405,193)(429,193){5}
input A;    //: /sn:0 {0}(353,155)(380,155)(380,154)(390,154){1}
//: {2}(394,154)(432,154){3}
//: {4}(392,156)(392,188)(429,188){5}
output C;    //: /sn:0 {0}(515,191)(450,191){1}
output S;    //: /sn:0 {0}(515,157)(453,157){1}
//: enddecls

  //: output g4 (C) @(512,191) /sn:0 /w:[ 0 ]
  //: input g3 (B) @(352,174) /sn:0 /w:[ 0 ]
  //: input g2 (A) @(351,155) /sn:0 /w:[ 0 ]
  xor g1 (.I0(A), .I1(B), .Z(S));   //: @(443,157) /sn:0 /delay:" 4" /w:[ 3 3 1 ]
  //: joint g6 (A) @(392, 154) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(405, 173) /w:[ 2 -1 1 4 ]
  //: output g5 (S) @(512,157) /sn:0 /w:[ 0 ]
  and g0 (.I0(A), .I1(B), .Z(C));   //: @(440,191) /sn:0 /delay:" 3" /w:[ 5 5 1 ]

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 {0}(197,204)(304,204)(304,213)(313,213){1}
wire w3;    //: /sn:0 /dp:1 {0}(498,267)(530,267){1}
wire w0;    //: /sn:0 {0}(197,250)(308,250)(308,258)(313,258){1}
wire w2;    //: /sn:0 {0}(498,240)(530,240){1}
//: enddecls

  led g4 (.I(w3));   //: @(537,267) /sn:0 /R:3 /w:[ 1 ] /type:0
  led g3 (.I(w2));   //: @(537,240) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: switch g2 (w0) @(180,250) /sn:0 /w:[ 0 ] /st:1
  Sumador_HA g1 (.B(w0), .A(w4), .C(w3), .S(w2));   //: @(314, 178) /sz:(183, 129) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: switch g0 (w4) @(180,204) /sn:0 /w:[ 0 ] /st:1

endmodule
