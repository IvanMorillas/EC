//: version "1.8.7"

module Sumador_HA(C, B, A, S);
//: interface  /sz:(183, 129) /bd:[ Li0>B(80/129) Li1>A(35/129) Ro0<C(89/129) Ro1<S(62/129) ]
input B;    //: /sn:0 {0}(354,174)(393,174)(393,173)(403,173){1}
//: {2}(407,173)(424,173)(424,159)(432,159){3}
//: {4}(405,175)(405,193)(429,193){5}
input A;    //: /sn:0 {0}(353,155)(380,155)(380,154)(390,154){1}
//: {2}(394,154)(432,154){3}
//: {4}(392,156)(392,188)(429,188){5}
output C;    //: /sn:0 {0}(515,191)(450,191){1}
output S;    //: /sn:0 {0}(515,157)(453,157){1}
//: enddecls

  //: output g4 (C) @(512,191) /sn:0 /w:[ 0 ]
  //: input g3 (B) @(352,174) /sn:0 /w:[ 0 ]
  //: input g2 (A) @(351,155) /sn:0 /w:[ 0 ]
  xor g1 (.I0(A), .I1(B), .Z(S));   //: @(443,157) /sn:0 /delay:" 4" /w:[ 3 3 1 ]
  //: joint g6 (A) @(392, 154) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(405, 173) /w:[ 2 -1 1 4 ]
  //: output g5 (S) @(512,157) /sn:0 /w:[ 0 ]
  and g0 (.I0(A), .I1(B), .Z(C));   //: @(440,191) /sn:0 /delay:" 3" /w:[ 5 5 1 ]

endmodule

module CPA(A, S, B, Cin);
//: interface  /sz:(40, 40) /bd:[ ]
input [3:0] B;    //: /sn:0 {0}(1157,146)(1089,146){1}
//: {2}(1088,146)(914,146){3}
//: {4}(913,146)(710,146){5}
//: {6}(709,146)(509,146){7}
//: {8}(508,146)(313,146){9}
input [3:0] A;    //: /sn:0 /dp:1 {0}(314,131)(469,131){1}
//: {2}(470,131)(696,131)(696,133){3}
//: {4}(696,134)(696,141)(879,141)(879,126)(894,126)(894,134){5}
//: {6}(894,135)(894,142)(965,142)(965,131)(1058,131){7}
//: {8}(1059,131)(1159,131){9}
input Cin;    //: /sn:0 {0}(1120,230)(1120,198)(1193,198){1}
output [4:0] S;    //: /sn:0 {0}(1397,420)(1250,420)(1250,425)(1240,425){1}
wire w16;    //: /sn:0 {0}(915,231)(915,158)(914,158)(914,150){1}
wire w13;    //: /sn:0 {0}(1106,339)(1106,360)(1006,360)(1006,213)(945,213)(945,231){1}
wire w6;    //: /sn:0 {0}(710,238)(710,150){1}
wire w7;    //: /sn:0 {0}(684,238)(684,134)(691,134){1}
wire w4;    //: /sn:0 {0}(479,329)(479,415)(1234,415){1}
wire w3;    //: /sn:0 {0}(526,329)(526,405)(1234,405){1}
wire w19;    //: /sn:0 {0}(887,333)(887,435)(1234,435){1}
wire w18;    //: /sn:0 {0}(930,333)(930,359)(838,359)(838,214)(756,214)(756,238){1}
wire w12;    //: /sn:0 {0}(1060,230)(1060,143)(1059,143)(1059,135){1}
wire w1;    //: /sn:0 {0}(509,237)(509,150){1}
wire w8;    //: /sn:0 {0}(739,330)(739,348)(625,348)(625,227)(543,227)(543,237){1}
wire w17;    //: /sn:0 {0}(881,231)(881,135)(889,135){1}
wire w14;    //: /sn:0 {0}(1066,339)(1066,445)(1234,445){1}
wire w11;    //: /sn:0 {0}(1091,230)(1091,158)(1089,158)(1089,150){1}
wire w2;    //: /sn:0 {0}(471,237)(471,143)(470,143)(470,135){1}
wire w9;    //: /sn:0 {0}(692,330)(692,425)(1234,425){1}
//: enddecls

  tran g8(.Z(w2), .I(A[3]));   //: @(470,129) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: input g4 (A) @(312,131) /sn:0 /w:[ 0 ]
  Sumador_FA g3 (.A(w17), .B(w16), .Cin(w13), .S(w19), .C(w18));   //: @(859, 232) /sz:(119, 100) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  //: output g16 (S) @(1394,420) /sn:0 /w:[ 0 ]
  Sumador_FA g2 (.A(w12), .B(w11), .Cin(Cin), .S(w14), .C(w13));   //: @(1040, 231) /sz:(110, 107) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Bo0<0 Bo1<0 ]
  Sumador_FA g1 (.A(w7), .B(w6), .Cin(w18), .S(w9), .C(w8));   //: @(660, 239) /sz:(132, 90) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  tran g10(.Z(w11), .I(B[0]));   //: @(1089,144) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g6(.Z(w17), .I(A[1]));   //: @(892,135) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:0
  //: input g9 (B) @(311,146) /sn:0 /w:[ 9 ]
  tran g7(.Z(w7), .I(A[2]));   //: @(694,134) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:0
  tran g12(.Z(w6), .I(B[2]));   //: @(710,144) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: input g14 (Cin) @(1195,198) /sn:0 /R:2 /w:[ 1 ]
  tran g11(.Z(w16), .I(B[1]));   //: @(914,144) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g5(.Z(w12), .I(A[0]));   //: @(1059,129) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  Sumador_FA g0 (.A(w2), .B(w1), .Cin(w8), .S(w4), .C(w3));   //: @(447, 238) /sz:(133, 90) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  concat g15 (.I0(w14), .I1(w19), .I2(w9), .I3(w4), .I4(w3), .Z(S));   //: @(1239,425) /sn:0 /w:[ 1 1 1 1 1 1 ] /dr:0
  tran g13(.Z(w1), .I(B[3]));   //: @(509,144) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1

endmodule

module Sumador_FA(B, A, C, S, Cin);
//: interface  /sz:(90, 70) /bd:[ Li0>Cin(51/70) Li1>B(33/70) Li2>A(13/70) Ro0<C(42/70) Ro1<S(17/70) ]
input B;    //: /sn:0 {0}(67,222)(120,222)(120,219)(130,219){1}
input A;    //: /sn:0 /dp:1 {0}(69,193)(120,193)(120,194)(130,194){1}
input Cin;    //: /sn:0 {0}(71,286)(327,286)(327,261)(337,261){1}
output C;    //: /sn:0 {0}(574,310)(544,310)(544,309)(514,309){1}
output S;    //: /sn:0 /dp:1 {0}(443,251)(584,251)(584,253)(594,253){1}
wire w7;    //: /sn:0 {0}(443,266)(483,266)(483,306)(493,306){1}
wire w2;    //: /sn:0 {0}(213,209)(273,209)(273,236)(337,236){1}
wire w9;    //: /sn:0 /dp:1 {0}(493,311)(264,311)(264,224)(213,224){1}
//: enddecls

  //: input g4 (B) @(65,222) /sn:0 /w:[ 0 ]
  //: input g3 (A) @(67,193) /sn:0 /w:[ 0 ]
  or g2 (.I0(w7), .I1(w9), .Z(C));   //: @(504,309) /sn:0 /delay:" 3" /w:[ 1 0 1 ]
  Sumador_HA g1 (.B(Cin), .A(w2), .C(w7), .S(S));   //: @(338, 218) /sz:(104, 70) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: output g6 (C) @(571,310) /sn:0 /w:[ 0 ]
  //: output g7 (S) @(591,253) /sn:0 /w:[ 1 ]
  //: input g5 (Cin) @(69,286) /sn:0 /w:[ 0 ]
  Sumador_HA g0 (.B(B), .A(A), .C(w9), .S(w2));   //: @(131, 176) /sz:(81, 70) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]

endmodule

module main;    //: root_module
wire [4:0] w4;    //: /sn:0 /dp:1 {0}(908,133)(908,213)(666,213){1}
wire [3:0] w0;    //: /sn:0 /dp:1 {0}(131,230)(131,243)(405,243){1}
wire w3;    //: /sn:0 {0}(216,289)(405,289){1}
wire [3:0] w2;    //: /sn:0 /dp:1 {0}(151,160)(151,184)(405,184){1}
//: enddecls

  //: dip g4 (w0) @(131,220) /sn:0 /w:[ 0 ] /st:6
  //: dip g3 (w2) @(151,150) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w3) @(199,289) /sn:0 /w:[ 0 ] /st:0
  led g1 (.I(w4));   //: @(908,126) /sn:0 /w:[ 0 ] /type:3
  CPA g0 (.Cin(w3), .B(w0), .A(w2), .S(w4));   //: @(406, 158) /sz:(259, 161) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Ro0<1 ]

endmodule
