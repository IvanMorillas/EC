//: version "1.8.7"

module CLL(C0, P1, C4, C3, C2, P2, P0, G1, G2, PG, P3, G0, G3, C1, GG);
//: interface  /sz:(818, 145) /bd:[ Ti0>G0(712/818) Ti1>P0(762/818) Ti2>G1(489/818) Ti3>P1(535/818) Ti4>P2(321/818) Ti5>G2(277/818) Ti6>P3(106/818) Ti7>G3(60/818) Ri0>C0(79/145) To0<C1(641/818) To1<C2(426/818) To2<C3(208/818) Lo0<C4(73/145) Bo0<PG(556/818) Bo1<GG(604/818) ]
input G2;    //: /sn:0 {0}(738,450)(332,450){1}
//: {2}(330,448)(330,351){3}
//: {4}(332,349)(342,349)(342,348)(968,348){5}
//: {6}(330,347)(330,117){7}
//: {8}(330,452)(330,538)(615,538){9}
output GG;    //: /sn:0 /dp:1 {0}(1024,561)(1064,561)(1064,532)(1101,532){1}
input C0;    //: /sn:0 {0}(568,122)(568,174){1}
//: {2}(570,176)(580,176)(580,175)(744,175){3}
//: {4}(568,178)(568,191){5}
//: {6}(570,193)(661,193)(661,192)(746,192){7}
//: {8}(568,195)(568,263){9}
//: {10}(570,265)(580,265)(580,266)(748,266){11}
//: {12}(568,267)(568,356){13}
//: {14}(570,358)(580,358)(580,356)(742,356){15}
//: {16}(568,360)(568,401){17}
input P1;    //: /sn:0 {0}(748,276)(393,276)(393,277)(383,277){1}
//: {2}(381,275)(381,225){3}
//: {4}(383,223)(393,223)(393,224)(746,224){5}
//: {6}(381,221)(381,203){7}
//: {8}(383,201)(393,201)(393,202)(746,202){9}
//: {10}(381,199)(381,120){11}
//: {12}(381,279)(381,301){13}
//: {14}(383,303)(393,303)(393,301)(748,301){15}
//: {16}(381,305)(381,363){17}
//: {18}(383,365)(393,365)(393,366)(742,366){19}
//: {20}(381,367)(381,390){21}
//: {22}(383,392)(741,392){23}
//: {24}(381,394)(381,465){25}
//: {26}(383,467)(412,467)(412,610)(845,610){27}
//: {28}(381,469)(381,490)(983,490){29}
output C3;    //: /sn:0 {0}(1153,349)(999,349)(999,340)(989,340){1}
output PG;    //: /sn:0 {0}(1129,479)(1046,479)(1046,485)(1069,485)(1069,492)(1004,492){1}
input G0;    //: /sn:0 {0}(520,121)(520,164){1}
//: {2}(522,166)(532,166)(532,155)(844,155){3}
//: {4}(520,168)(520,219){5}
//: {6}(522,221)(532,221)(532,219)(746,219){7}
//: {8}(520,223)(520,293){9}
//: {10}(522,295)(532,295)(532,296)(748,296){11}
//: {12}(520,297)(520,387)(523,387){13}
//: {14}(527,387)(741,387){15}
//: {16}(525,389)(525,605)(845,605){17}
output C4;    //: /sn:0 /dp:1 {0}(974,375)(1148,375)(1148,413)(1158,413){1}
output C2;    //: /sn:0 /dp:1 {0}(964,230)(1105,230)(1105,297)(1153,297){1}
input P3;    //: /sn:0 {0}(650,529)(232,529){1}
//: {2}(230,527)(230,471){3}
//: {4}(232,469)(241,469)(241,442)(232,442){5}
//: {6}(230,440)(230,427){7}
//: {8}(232,425)(739,425){9}
//: {10}(230,423)(230,404){11}
//: {12}(232,402)(741,402){13}
//: {14}(230,400)(230,378){15}
//: {16}(232,376)(742,376){17}
//: {18}(230,374)(230,120){19}
//: {20}(228,442)(218,442)(218,500)(983,500){21}
//: {22}(230,444)(230,445)(738,445){23}
//: {24}(230,467)(230,457)(245,457)(245,620)(845,620){25}
//: {26}(230,531)(230,543)(615,543){27}
input G1;    //: /sn:0 {0}(739,415)(434,415){1}
//: {2}(430,415)(427,415)(427,333){3}
//: {4}(429,331)(439,331)(439,330)(746,330){5}
//: {6}(427,329)(427,237){7}
//: {8}(429,235)(943,235){9}
//: {10}(427,233)(427,119){11}
//: {12}(432,417)(432,519)(650,519){13}
input G3;    //: /sn:0 {0}(1003,569)(255,569)(255,455){1}
//: {2}(257,453)(945,453)(945,385)(953,385){3}
//: {4}(255,451)(255,122){5}
input P0;    //: /sn:0 {0}(983,485)(475,485)(475,361){1}
//: {2}(477,359)(487,359)(487,361)(742,361){3}
//: {4}(475,357)(475,270){5}
//: {6}(477,268)(487,268)(487,271)(748,271){7}
//: {8}(475,266)(475,199){9}
//: {10}(477,197)(746,197){11}
//: {12}(475,195)(475,173){13}
//: {14}(477,171)(487,171)(487,170)(744,170){15}
//: {16}(475,169)(475,120){17}
output C1;    //: /sn:0 /dp:1 {0}(865,158)(1142,158)(1142,236)(1157,236){1}
input P2;    //: /sn:0 {0}(845,615)(306,615)(306,519)(297,519){1}
//: {2}(295,517)(295,482)(287,482){3}
//: {4}(285,480)(285,422){5}
//: {6}(287,420)(739,420){7}
//: {8}(285,418)(285,399){9}
//: {10}(287,397)(741,397){11}
//: {12}(285,395)(285,372){13}
//: {14}(287,370)(297,370)(297,371)(742,371){15}
//: {16}(285,368)(285,339){17}
//: {18}(287,337)(297,337)(297,335)(746,335){19}
//: {20}(285,335)(285,309){21}
//: {22}(287,307)(297,307)(297,306)(748,306){23}
//: {24}(285,305)(285,285){25}
//: {26}(287,283)(297,283)(297,281)(748,281){27}
//: {28}(285,281)(285,121){29}
//: {30}(285,484)(285,495)(983,495){31}
//: {32}(295,521)(295,524)(650,524){33}
wire w16;    //: /sn:0 {0}(671,524)(690,524)(690,559)(1003,559){1}
wire w13;    //: /sn:0 {0}(762,394)(772,394)(772,370)(953,370){1}
wire w7;    //: /sn:0 {0}(763,366)(943,366)(943,365)(953,365){1}
wire w3;    //: /sn:0 {0}(767,197)(933,197)(933,225)(943,225){1}
wire w20;    //: /sn:0 {0}(759,448)(788,448)(788,380)(953,380){1}
wire w12;    //: /sn:0 {0}(769,301)(928,301)(928,338)(968,338){1}
wire w10;    //: /sn:0 {0}(767,222)(889,222)(889,230)(943,230){1}
wire w21;    //: /sn:0 {0}(636,541)(675,541)(675,564)(1003,564){1}
wire w1;    //: /sn:0 /dp:1 {0}(844,160)(828,160)(828,173)(765,173){1}
wire w8;    //: /sn:0 {0}(769,273)(958,273)(958,333)(968,333){1}
wire w17;    //: /sn:0 {0}(760,420)(777,420)(777,375)(953,375){1}
wire w15;    //: /sn:0 {0}(767,333)(913,333)(913,343)(968,343){1}
wire w9;    //: /sn:0 {0}(866,612)(992,612)(992,554)(1003,554){1}
//: enddecls

  //: input g4 (C0) @(568,120) /sn:0 /R:3 /w:[ 0 ]
  //: input g8 (P1) @(381,118) /sn:0 /R:3 /w:[ 11 ]
  and g44 (.I0(G1), .I1(P2), .I2(P3), .Z(w17));   //: @(750,420) /sn:0 /delay:" 3" /w:[ 0 7 9 0 ]
  //: output g3 (C4) @(1155,413) /sn:0 /w:[ 1 ]
  or g16 (.I0(G0), .I1(w1), .Z(C1));   //: @(855,158) /sn:0 /delay:" 3" /w:[ 3 0 0 ]
  //: joint g47 (P0) @(475, 359) /w:[ 2 4 -1 1 ]
  //: joint g17 (G0) @(520, 166) /w:[ 2 1 -1 4 ]
  //: joint g26 (G1) @(427, 235) /w:[ 8 10 -1 7 ]
  //: output g2 (C3) @(1150,349) /sn:0 /w:[ 0 ]
  //: joint g23 (P1) @(381, 201) /w:[ 8 10 -1 7 ]
  and g30 (.I0(G1), .I1(P2), .Z(w15));   //: @(757,333) /sn:0 /delay:" 3" /w:[ 5 19 0 ]
  //: output g1 (C2) @(1150,297) /sn:0 /w:[ 1 ]
  //: joint g24 (G0) @(520, 221) /w:[ 6 5 -1 8 ]
  //: joint g39 (P2) @(285, 337) /w:[ 18 20 -1 17 ]
  or g60 (.I0(w9), .I1(w16), .I2(w21), .I3(G3), .Z(GG));   //: @(1014,561) /sn:0 /delay:" 3" /w:[ 1 1 1 0 0 ]
  and g29 (.I0(G0), .I1(P1), .I2(P2), .Z(w12));   //: @(759,301) /sn:0 /delay:" 3" /w:[ 11 15 23 0 ]
  //: joint g51 (P3) @(230, 376) /w:[ 16 18 -1 15 ]
  //: joint g70 (P2) @(295, 519) /w:[ 1 2 -1 32 ]
  and g18 (.I0(C0), .I1(P0), .I2(P1), .Z(w3));   //: @(757,197) /sn:0 /delay:" 3" /w:[ 7 11 9 0 ]
  //: joint g65 (G2) @(330, 450) /w:[ 1 2 -1 8 ]
  //: input g10 (P2) @(285,119) /sn:0 /R:3 /w:[ 29 ]
  //: joint g25 (P1) @(381, 223) /w:[ 4 6 -1 3 ]
  and g64 (.I0(G2), .I1(P3), .Z(w21));   //: @(626,541) /sn:0 /w:[ 9 27 0 ]
  //: joint g72 (G0) @(525, 387) /w:[ 14 -1 13 16 ]
  //: joint g49 (P2) @(285, 370) /w:[ 14 16 -1 13 ]
  //: input g6 (P0) @(475,118) /sn:0 /R:3 /w:[ 17 ]
  //: joint g50 (P2) @(285, 397) /w:[ 10 12 -1 9 ]
  //: joint g68 (G1) @(432, 415) /w:[ 1 -1 2 12 ]
  //: joint g58 (P2) @(285, 420) /w:[ 6 8 -1 5 ]
  and g56 (.I0(P0), .I1(P1), .I2(P2), .I3(P3), .Z(PG));   //: @(994,492) /sn:0 /delay:" 3" /w:[ 0 29 31 21 1 ]
  //: input g7 (G1) @(427,117) /sn:0 /R:3 /w:[ 11 ]
  //: input g9 (G2) @(330,115) /sn:0 /R:3 /w:[ 7 ]
  //: joint g35 (G0) @(520, 295) /w:[ 10 9 -1 12 ]
  //: joint g71 (P1) @(381, 467) /w:[ 26 25 -1 28 ]
  //: joint g59 (P3) @(230, 442) /w:[ 5 6 20 22 ]
  //: joint g22 (P0) @(475, 197) /w:[ 10 12 -1 9 ]
  //: joint g31 (C0) @(568, 265) /w:[ 10 9 -1 12 ]
  //: joint g67 (P2) @(285, 482) /w:[ 3 4 -1 30 ]
  //: output g54 (PG) @(1126,479) /sn:0 /w:[ 0 ]
  //: joint g33 (P1) @(381, 277) /w:[ 1 2 -1 12 ]
  //: joint g36 (P1) @(381, 303) /w:[ 14 13 -1 16 ]
  or g41 (.I0(w7), .I1(w13), .I2(w17), .I3(w20), .I4(G3), .Z(C4));   //: @(964,375) /sn:0 /delay:" 3" /w:[ 1 1 1 1 3 0 ]
  and g45 (.I0(P3), .I1(G2), .Z(w20));   //: @(749,448) /sn:0 /delay:" 3" /w:[ 23 0 0 ]
  //: joint g69 (P3) @(230, 529) /w:[ 1 2 -1 26 ]
  //: joint g40 (G2) @(330, 349) /w:[ 4 6 -1 3 ]
  and g42 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .I4(P3), .Z(w7));   //: @(753,366) /sn:0 /delay:" 3" /w:[ 15 3 19 15 17 0 ]
  //: joint g52 (P3) @(230, 402) /w:[ 12 14 -1 11 ]
  //: joint g66 (P3) @(230, 469) /w:[ 4 24 -1 3 ]
  //: input g12 (P3) @(230,118) /sn:0 /R:3 /w:[ 19 ]
  //: joint g57 (P1) @(381, 392) /w:[ 22 21 -1 24 ]
  and g28 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .Z(w8));   //: @(759,273) /sn:0 /delay:" 3" /w:[ 11 7 0 27 0 ]
  //: joint g34 (P2) @(285, 283) /w:[ 26 28 -1 25 ]
  //: joint g46 (C0) @(568, 358) /w:[ 14 13 -1 16 ]
  //: input g5 (G0) @(520,119) /sn:0 /R:3 /w:[ 0 ]
  //: input g11 (G3) @(255,120) /sn:0 /R:3 /w:[ 5 ]
  //: joint g14 (P0) @(475, 171) /w:[ 14 16 -1 13 ]
  //: joint g61 (G3) @(255, 453) /w:[ 2 4 -1 1 ]
  or g19 (.I0(w3), .I1(w10), .I2(G1), .Z(C2));   //: @(954,230) /sn:0 /delay:" 3" /w:[ 1 1 9 0 ]
  //: joint g21 (C0) @(568, 193) /w:[ 6 5 -1 8 ]
  and g20 (.I0(G0), .I1(P1), .Z(w10));   //: @(757,222) /sn:0 /delay:" 3" /w:[ 7 5 0 ]
  //: joint g32 (P0) @(475, 268) /w:[ 6 8 -1 5 ]
  and g63 (.I0(G1), .I1(P2), .I2(P3), .Z(w16));   //: @(661,524) /sn:0 /w:[ 13 33 0 0 ]
  //: joint g15 (C0) @(568, 176) /w:[ 2 1 -1 4 ]
  //: output g0 (C1) @(1154,236) /sn:0 /w:[ 1 ]
  //: joint g38 (G1) @(427, 331) /w:[ 4 6 -1 3 ]
  and g43 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w13));   //: @(752,394) /sn:0 /delay:" 3" /w:[ 15 23 11 13 0 ]
  or g27 (.I0(w8), .I1(w12), .I2(w15), .I3(G2), .Z(C3));   //: @(979,340) /sn:0 /delay:" 3" /w:[ 1 1 1 5 1 ]
  //: joint g48 (P1) @(381, 365) /w:[ 18 17 -1 20 ]
  and g62 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w9));   //: @(856,612) /sn:0 /w:[ 17 27 0 25 0 ]
  //: joint g37 (P2) @(285, 307) /w:[ 22 24 -1 21 ]
  //: output g55 (GG) @(1098,532) /sn:0 /w:[ 1 ]
  and g13 (.I0(P0), .I1(C0), .Z(w1));   //: @(755,173) /sn:0 /delay:" 3" /w:[ 15 3 1 ]
  //: joint g53 (P3) @(230, 425) /w:[ 8 10 -1 7 ]

endmodule

module PFA(Pi, Cin, B, S, Gi, A);
//: interface  /sz:(181, 159) /bd:[ Ti0>Cin(44/181) Ti1>B(106/181) Ti2>A(134/181) Bo0<Gi(49/181) Bo1<Pi(98/181) Bo2<S(129/181) ]
input B;    //: /sn:0 {0}(524,190)(573,190){1}
//: {2}(577,190)(698,190)(698,182)(708,182){3}
//: {4}(575,192)(575,273){5}
//: {6}(577,275)(688,275)(688,260)(800,260){7}
//: {8}(575,277)(575,288)(798,288){9}
output Gi;    //: /sn:0 /dp:1 {0}(819,291)(933,291){1}
input A;    //: /sn:0 {0}(526,152)(593,152){1}
//: {2}(597,152)(698,152)(698,177)(708,177){3}
//: {4}(595,154)(595,247){5}
//: {6}(597,249)(790,249)(790,255)(800,255){7}
//: {8}(595,251)(595,293)(798,293){9}
input Cin;    //: /sn:0 {0}(529,233)(770,233)(770,208)(802,208){1}
output Pi;    //: /sn:0 {0}(930,258)(821,258){1}
output S;    //: /sn:0 /dp:1 {0}(823,206)(930,206){1}
wire w2;    //: /sn:0 {0}(729,180)(792,180)(792,203)(802,203){1}
//: enddecls

  xor g4 (.I0(w2), .I1(Cin), .Z(S));   //: @(813,206) /sn:0 /delay:" 4" /w:[ 1 1 0 ]
  //: output g8 (Pi) @(927,258) /sn:0 /w:[ 0 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(719,180) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: input g2 (Cin) @(527,233) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(522,190) /sn:0 /w:[ 0 ]
  //: joint g10 (A) @(595, 152) /w:[ 2 -1 1 4 ]
  or g6 (.I0(A), .I1(B), .Z(Pi));   //: @(811,258) /sn:0 /delay:" 3" /w:[ 7 7 1 ]
  //: output g7 (S) @(927,206) /sn:0 /w:[ 1 ]
  //: output g9 (Gi) @(930,291) /sn:0 /w:[ 1 ]
  //: joint g12 (A) @(595, 249) /w:[ 6 5 -1 8 ]
  and g5 (.I0(B), .I1(A), .Z(Gi));   //: @(809,291) /sn:0 /delay:" 3" /w:[ 9 9 0 ]
  //: joint g11 (B) @(575, 190) /w:[ 2 -1 1 4 ]
  //: input g0 (A) @(524,152) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(575, 275) /w:[ 6 5 -1 8 ]

endmodule

module CLA_16(Cin, PG, Cout, S, A, GG, B);
//: interface  /sz:(224, 223) /bd:[ Ti0>A[15:0](179/224) Ti1>B[15:0](134/224) Ti2>Cin(67/224) Bo0<S[15:0](174/224) Bo1<Cout(144/224) Bo2<PG(42/224) Bo3<GG(85/224) ]
input [15:0] B;    //: /sn:0 {0}(1003,-210)(849,-210){1}
//: {2}(848,-210)(530,-210){3}
//: {4}(529,-210)(223,-210)(223,-214){5}
//: {6}(223,-215)(223,-230)(-9,-230)(-9,-210)(-97,-210){7}
//: {8}(-98,-210)(-261,-210){9}
output GG;    //: /sn:0 /dp:1 {0}(699,592)(699,648)(717,648){1}
input [15:0] A;    //: /sn:0 /dp:3 {0}(-263,-251)(2,-251){1}
//: {2}(3,-251)(311,-251){3}
//: {4}(312,-251)(620,-251)(620,-255){5}
//: {6}(620,-256)(620,-260)(778,-260)(778,-251)(950,-251){7}
//: {8}(951,-251)(1003,-251){9}
output PG;    //: /sn:0 {0}(658,647)(634,647)(634,592){1}
input Cin;    //: /sn:0 {0}(1108,125)(1108,129)(1081,129){1}
//: {2}(1077,129)(1041,129){3}
//: {4}(1079,131)(1079,503)(990,503){5}
output Cout;    //: /sn:0 {0}(-236,504)(-236,495)(-120,495){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(1137,358)(1196,358)(1196,357)(1270,357){1}
wire [3:0] w16;    //: /sn:0 {0}(1131,343)(14,343)(14,280){1}
wire [3:0] w13;    //: /sn:0 /dp:1 {0}(1131,353)(322,353)(322,282){1}
wire [3:0] w6;    //: /sn:0 {0}(633,96)(633,-255)(624,-255){1}
wire [3:0] w7;    //: /sn:0 {0}(530,96)(530,-206){1}
wire w25;    //: /sn:0 {0}(221,282)(221,339)(224,339)(224,398){1}
wire [3:0] w3;    //: /sn:0 {0}(312,87)(312,-247){1}
wire [3:0] w0;    //: /sn:0 {0}(951,95)(951,-247){1}
wire w30;    //: /sn:0 {0}(-36,280)(-36,391)(-44,391)(-44,398){1}
wire [3:0] w10;    //: /sn:0 /dp:1 {0}(1131,373)(961,373)(961,290){1}
wire w23;    //: /sn:0 {0}(272,282)(272,342)(281,342)(281,398){1}
wire w24;    //: /sn:0 {0}(542,291)(542,355)(554,355)(554,398){1}
wire w31;    //: /sn:0 {0}(-87,280)(-87,391)(-86,391)(-86,398){1}
wire [3:0] w1;    //: /sn:0 {0}(848,95)(848,-198)(849,-198)(849,-206){1}
wire [3:0] w8;    //: /sn:0 {0}(209,87)(209,-214)(218,-214){1}
wire [3:0] w27;    //: /sn:0 {0}(-99,85)(-99,-198)(-97,-198)(-97,-206){1}
wire w17;    //: /sn:0 {0}(98,398)(98,119)(94,119){1}
wire w14;    //: /sn:0 {0}(723,130)(767,130)(767,398){1}
wire [3:0] w11;    //: /sn:0 {0}(1131,363)(643,363)(643,291){1}
wire w2;    //: /sn:0 /dp:1 {0}(911,290)(911,351)(913,351)(913,398){1}
wire w15;    //: /sn:0 /dp:1 {0}(402,121)(418,121)(418,398){1}
wire w5;    //: /sn:0 {0}(860,290)(860,356)(845,356)(845,398){1}
wire [3:0] w26;    //: /sn:0 {0}(4,85)(4,-239)(3,-239)(3,-247){1}
wire w9;    //: /sn:0 {0}(604,398)(604,348)(593,348)(593,291){1}
//: enddecls

  concat g8 (.I0(w10), .I1(w11), .I2(w13), .I3(w16), .Z(S));   //: @(1136,358) /sn:0 /w:[ 0 0 0 0 0 ] /dr:0
  //: input g4 (Cin) @(1108,123) /sn:0 /R:3 /w:[ 0 ]
  tran g16(.Z(w6), .I(A[7:4]));   //: @(618,-255) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:1
  CLA g3 (.B(w7), .A(w6), .Cin(w14), .GG(w24), .PG(w9), .S(w11));   //: @(454, 97) /sz:(268, 193) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<0 Bo1<1 Bo2<1 ]
  tran g17(.Z(w3), .I(A[11:8]));   //: @(312,-253) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: joint g2 (Cin) @(1079, 129) /w:[ 1 -1 2 4 ]
  CLL g1 (.G3(w31), .P3(w30), .G2(w25), .P2(w23), .P1(w9), .G1(w24), .P0(w2), .G0(w5), .C0(Cin), .C3(w17), .C2(w15), .C1(w14), .C4(Cout), .GG(GG), .PG(PG));   //: @(-119, 399) /sz:(1108, 192) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>0 Ti5>1 Ti6>1 Ti7>1 Ri0>5 To0<0 To1<1 To2<1 Lo0<1 Bo0<0 Bo1<1 ]
  tran g18(.Z(w1), .I(B[3:0]));   //: @(849,-212) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  //: output g10 (PG) @(655,647) /sn:0 /w:[ 0 ]
  CLA g6 (.B(w27), .A(w26), .Cin(w17), .GG(w31), .PG(w30), .S(w16));   //: @(-175, 86) /sz:(268, 193) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<1 ]
  //: output g9 (Cout) @(-236,501) /sn:0 /R:3 /w:[ 0 ]
  //: output g7 (S) @(1267,357) /sn:0 /w:[ 1 ]
  //: input g12 (A) @(-265,-251) /sn:0 /w:[ 0 ]
  tran g14(.Z(w0), .I(A[3:0]));   //: @(951,-253) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: output g11 (GG) @(714,648) /sn:0 /w:[ 1 ]
  CLA g5 (.B(w8), .A(w3), .Cin(w15), .GG(w25), .PG(w23), .S(w13));   //: @(133, 88) /sz:(268, 193) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Bo0<0 Bo1<0 Bo2<1 ]
  tran g21(.Z(w27), .I(B[15:12]));   //: @(-97,-212) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  tran g19(.Z(w7), .I(B[7:4]));   //: @(530,-212) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g20(.Z(w8), .I(B[11:8]));   //: @(221,-214) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:0
  tran g15(.Z(w26), .I(A[15:12]));   //: @(3,-253) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  CLA g0 (.B(w1), .A(w0), .Cin(Cin), .GG(w5), .PG(w2), .S(w10));   //: @(772, 96) /sz:(268, 193) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>3 Bo0<0 Bo1<0 Bo2<1 ]
  //: input g13 (B) @(-263,-210) /sn:0 /w:[ 9 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(731,464)(731,500){1}
wire [15:0] w7;    //: /sn:0 {0}(867,211)(867,225)(825,225)(825,239){1}
wire w4;    //: /sn:0 {0}(790,464)(790,501){1}
wire [15:0] w0;    //: /sn:0 /dp:1 {0}(779,215)(779,230)(780,230)(780,239){1}
wire w1;    //: /sn:0 {0}(648,190)(713,190)(713,239){1}
wire [15:0] w2;    //: /sn:0 {0}(967,482)(967,492)(820,492)(820,464){1}
wire w5;    //: /sn:0 {0}(688,464)(688,501){1}
//: enddecls

  led g4 (.I(w2));   //: @(967,475) /sn:0 /w:[ 0 ] /type:3
  //: switch g3 (w1) @(631,190) /sn:0 /w:[ 0 ] /st:0
  //: dip g2 (w0) @(779,205) /sn:0 /w:[ 0 ] /st:0
  //: dip g1 (w7) @(867,201) /sn:0 /w:[ 0 ] /st:0
  led g6 (.I(w6));   //: @(731,507) /sn:0 /R:2 /w:[ 1 ] /type:0
  led g7 (.I(w5));   //: @(688,508) /sn:0 /R:2 /w:[ 1 ] /type:0
  led g5 (.I(w4));   //: @(790,508) /sn:0 /R:2 /w:[ 1 ] /type:0
  CLA_16 g0 (.Cin(w1), .B(w0), .A(w7), .GG(w6), .PG(w5), .Cout(w4), .S(w2));   //: @(646, 240) /sz:(224, 223) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Bo0<0 Bo1<0 Bo2<0 Bo3<1 ]

endmodule

module CLA(A, S, Cout, Cin, GG, PG, B);
//: interface  /sz:(268, 193) /bd:[ Ti0>A[3:0](179/268) Ti1>B[3:0](76/268) Ri0>Cin(33/193) Bo0<S[3:0](189/268) Bo1<PG(139/268) Bo2<GG(88/268) ]
input [3:0] B;    //: /sn:0 {0}(-161,-173)(-109,-173){1}
//: {2}(-108,-173)(116,-173){3}
//: {4}(117,-173)(330,-173){5}
//: {6}(331,-173)(542,-173){7}
//: {8}(543,-173)(654,-173){9}
output GG;    //: /sn:0 {0}(388,489)(388,540){1}
input [3:0] A;    //: /sn:0 {0}(-159,-203)(-82,-203){1}
//: {2}(-81,-203)(143,-203){3}
//: {4}(144,-203)(252,-203)(252,-202)(359,-202){5}
//: {6}(360,-202)(465,-202)(465,-203)(568,-203){7}
//: {8}(569,-203)(650,-203){9}
output PG;    //: /sn:0 {0}(340,489)(340,542){1}
input Cin;    //: /sn:0 /dp:1 {0}(481,48)(481,27)(737,27){1}
//: {2}(741,27)(841,27){3}
//: {4}(739,29)(739,422)(603,422){5}
output Cout;    //: /sn:0 {0}(-263,414)(-228,414)(-228,416)(-217,416){1}
output [3:0] S;    //: /sn:0 {0}(696,272)(666,272)(666,262)(636,262){1}
wire w16;    //: /sn:0 {0}(105,212)(105,342){1}
wire w13;    //: /sn:0 {0}(117,51)(117,-169){1}
wire w7;    //: /sn:0 {0}(331,45)(331,-169){1}
wire w22;    //: /sn:0 {0}(-117,213)(-117,332)(-110,332)(-110,342){1}
wire w36;    //: /sn:0 /dp:1 {0}(269,45)(269,37)(425,37)(425,342){1}
wire w0;    //: /sn:0 /dp:1 {0}(210,342)(210,43)(55,43)(55,51){1}
wire w3;    //: /sn:0 {0}(486,209)(486,332)(496,332)(496,342){1}
wire w20;    //: /sn:0 {0}(-81,52)(-81,-199){1}
wire w19;    //: /sn:0 {0}(-109,52)(-109,-161)(-108,-161)(-108,-169){1}
wire w12;    //: /sn:0 /dp:1 {0}(-8,342)(-8,44)(-171,44)(-171,52){1}
wire w23;    //: /sn:0 {0}(-86,213)(-86,247)(630,247){1}
wire w10;    //: /sn:0 {0}(323,206)(323,331)(319,331)(319,342){1}
wire w21;    //: /sn:0 {0}(-166,213)(-166,332)(-156,332)(-156,342){1}
wire w1;    //: /sn:0 {0}(543,48)(543,-169){1}
wire w8;    //: /sn:0 /dp:1 {0}(359,45)(359,-196)(360,-196)(360,-198){1}
wire w17;    //: /sn:0 {0}(140,212)(140,257)(630,257){1}
wire w14;    //: /sn:0 {0}(145,51)(145,-191)(144,-191)(144,-199){1}
wire w11;    //: /sn:0 {0}(354,206)(354,267)(630,267){1}
wire w2;    //: /sn:0 {0}(571,48)(571,-191)(569,-191)(569,-199){1}
wire w15;    //: /sn:0 {0}(60,212)(60,332)(61,332)(61,342){1}
wire w5;    //: /sn:0 {0}(566,209)(566,277)(630,277){1}
wire w26;    //: /sn:0 /dp:1 {0}(546,342)(546,332)(535,332)(535,209){1}
wire w9;    //: /sn:0 {0}(274,206)(274,332)(273,332)(273,342){1}
//: enddecls

  //: input g8 (A) @(-161,-203) /sn:0 /w:[ 0 ]
  CLL g4 (.G3(w21), .P3(w22), .G2(w15), .P2(w16), .P1(w10), .G1(w9), .P0(w26), .G0(w3), .C0(Cin), .C3(w12), .C2(w0), .C1(w36), .C4(Cout), .GG(GG), .PG(PG));   //: @(-216, 343) /sz:(818, 145) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>0 Ti7>1 Ri0>5 To0<0 To1<0 To2<1 Lo0<1 Bo0<0 Bo1<0 ]
  tran g16(.Z(w19), .I(B[3]));   //: @(-108,-175) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  PFA g3 (.A(w20), .B(w19), .Cin(w12), .S(w23), .Pi(w22), .Gi(w21));   //: @(-215, 53) /sz:(181, 159) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 Bo2<0 ]
  tran g17(.Z(w7), .I(B[1]));   //: @(331,-175) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  PFA g2 (.A(w14), .B(w13), .Cin(w0), .S(w17), .Pi(w16), .Gi(w15));   //: @(11, 52) /sz:(181, 159) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 Bo2<0 ]
  PFA g1 (.A(w8), .B(w7), .Cin(w36), .S(w11), .Pi(w10), .Gi(w9));   //: @(226, 46) /sz:(180, 159) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  //: output g18 (S) @(693,272) /sn:0 /w:[ 0 ]
  tran g10(.Z(w14), .I(A[2]));   //: @(144,-205) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: joint g6 (Cin) @(739, 27) /w:[ 2 -1 1 4 ]
  tran g9(.Z(w2), .I(A[0]));   //: @(569,-205) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: output g7 (Cout) @(-260,414) /sn:0 /R:2 /w:[ 0 ]
  tran g12(.Z(w8), .I(A[1]));   //: @(360,-204) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g14(.Z(w1), .I(B[0]));   //: @(543,-175) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g11(.Z(w20), .I(A[3]));   //: @(-81,-205) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: input g5 (Cin) @(843,27) /sn:0 /R:2 /w:[ 3 ]
  //: output g21 (GG) @(388,537) /sn:0 /R:3 /w:[ 1 ]
  concat g19 (.I0(w5), .I1(w11), .I2(w17), .I3(w23), .Z(S));   //: @(635,262) /sn:0 /w:[ 1 1 1 1 1 ] /dr:0
  //: output g20 (PG) @(340,539) /sn:0 /R:3 /w:[ 1 ]
  tran g15(.Z(w13), .I(B[2]));   //: @(117,-175) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  PFA g0 (.A(w2), .B(w1), .Cin(Cin), .S(w5), .Pi(w26), .Gi(w3));   //: @(437, 49) /sz:(181, 159) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Bo0<0 Bo1<1 Bo2<0 ]
  //: input g13 (B) @(-163,-173) /sn:0 /w:[ 0 ]

endmodule
