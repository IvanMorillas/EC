//: version "1.8.7"

module MEM(WriteData, MemRead, ReadData, MemWrite, Address);
//: interface  /sz:(102, 199) /bd:[ Ti0>MemWrite(55/102) Li0>WriteData[31:0](166/199) Li1>Address[31:0](70/199) Bi0>MemRead(54/102) Ro0<ReadData[31:0](96/199) ]
output [31:0] ReadData;    //: /sn:0 /dp:1 {0}(483,166)(483,235){1}
//: {2}(485,237)(647,237){3}
//: {4}(481,237)(390,237){5}
input [31:0] WriteData;    //: /sn:0 {0}(369,81)(483,81)(483,150){1}
supply0 w3;    //: /sn:0 {0}(398,361)(398,349)(382,349)(382,339){1}
input MemWrite;    //: /sn:0 {0}(201,134)(272,134){1}
supply0 w1;    //: /sn:0 {0}(366,283)(366,264){1}
supply0 w2;    //: /sn:0 {0}(241,114)(252,114)(252,129)(272,129){1}
input MemRead;    //: /sn:0 {0}(377,384)(377,339){1}
input [31:0] Address;    //: /sn:0 {0}(199,239)(355,239){1}
wire w6;    //: /sn:0 {0}(380,318)(380,264){1}
wire w7;    //: /sn:0 {0}(293,132)(371,132){1}
//: {2}(375,132)(498,132)(498,158)(488,158){3}
//: {4}(373,134)(373,146){5}
wire w9;    //: /sn:0 {0}(373,162)(373,214){1}
//: enddecls

  //: input g4 (WriteData) @(367,81) /sn:0 /w:[ 0 ]
  //: joint g8 (ReadData) @(483, 237) /w:[ 2 1 4 -1 ]
  //: input g3 (MemRead) @(377,386) /sn:0 /R:1 /w:[ 0 ]
  //: output g2 (ReadData) @(644,237) /sn:0 /w:[ 3 ]
  //: input g1 (MemWrite) @(199,134) /sn:0 /w:[ 0 ]
  not g10 (.I(w7), .Z(w9));   //: @(373,152) /sn:0 /R:3 /w:[ 5 0 ]
  //: supply0 g6 (w1) @(366,289) /sn:0 /w:[ 0 ]
  bufif1 g7 (.Z(ReadData), .I(WriteData), .E(w7));   //: @(483,156) /sn:0 /R:3 /w:[ 0 1 3 ]
  and g9 (.I0(w2), .I1(MemWrite), .Z(w7));   //: @(283,132) /sn:0 /w:[ 1 1 0 ]
  //: supply0 g12 (w2) @(235,114) /sn:0 /R:3 /w:[ 0 ]
  ram g5 (.A(Address), .D(ReadData), .WE(w9), .OE(w6), .CS(w1));   //: @(373,238) /sn:0 /w:[ 1 5 1 1 1 ]
  //: joint g11 (w7) @(373, 132) /w:[ 2 -1 1 4 ]
  //: supply0 g14 (w3) @(398,367) /sn:0 /w:[ 0 ]
  //: input g0 (Address) @(197,239) /sn:0 /w:[ 0 ]
  nand g13 (.I0(MemRead), .I1(w3), .Z(w6));   //: @(380,328) /sn:0 /R:1 /w:[ 1 1 0 ]

endmodule

module READ(RegDst, Data1, RegMux, Reg2, Reg1, clk, Data, Data2, clr, RegWrite, ESignExt, SSignExt);
//: interface  /sz:(244, 247) /bd:[ Ti0>clr(131/244) Ti1>clr(131/244) Li0>Reg1[4:0](31/247) Li1>Reg2[4:0](77/247) Li2>RegMux[4:0](117/247) Li3>RegDst(152/247) Li4>ESignExt[15:0](202/247) Li5>ESignExt[15:0](202/247) Li6>RegDst(152/247) Li7>RegMux[4:0](117/247) Li8>Reg2[4:0](77/247) Li9>Reg1[4:0](31/247) Bi0>Data[31:0](62/244) Bi1>clk(160/244) Bi2>RegWrite(116/244) Bi3>RegWrite(116/244) Bi4>clk(160/244) Bi5>Data[31:0](62/244) Ro0<Data1[31:0](63/247) Ro1<Data2[31:0](126/247) Ro2<SSignExt[31:0](196/247) Ro3<SSignExt[31:0](196/247) Ro4<Data2[31:0](126/247) Ro5<Data1[31:0](63/247) ]
output [31:0] Data2;    //: /sn:0 {0}(885,395)(779,395){1}
input [4:0] Reg1;    //: /sn:0 {0}(366,288)(630,288){1}
output [31:0] SSignExt;    //: /sn:0 /dp:1 {0}(752,613)(825,613){1}
input [4:0] RegMux;    //: /sn:0 {0}(371,374)(472,374){1}
output [31:0] Data1;    //: /sn:0 {0}(887,303)(779,303){1}
input RegDst;    //: /sn:0 {0}(367,419)(488,419)(488,387){1}
input [4:0] Reg2;    //: /sn:0 {0}(368,328)(452,328){1}
//: {2}(456,328)(630,328){3}
//: {4}(454,330)(454,354)(472,354){5}
input RegWrite;    //: /sn:0 {0}(671,504)(671,439){1}
input clr;    //: /sn:0 {0}(687,170)(697,170)(697,255){1}
input clk;    //: /sn:0 {0}(739,505)(739,439){1}
input [31:0] Data;    //: /sn:0 {0}(565,404)(630,404){1}
input [15:0] ESignExt;    //: /sn:0 {0}(604,614)(657,614){1}
wire [4:0] w12;    //: /sn:0 {0}(501,364)(630,364){1}
//: enddecls

  //: input g4 (RegDst) @(365,419) /sn:0 /w:[ 0 ]
  //: output g8 (Data1) @(884,303) /sn:0 /w:[ 0 ]
  //: input g3 (RegMux) @(369,374) /sn:0 /w:[ 0 ]
  //: input g2 (Reg2) @(366,328) /sn:0 /w:[ 0 ]
  //: input g1 (Reg1) @(364,288) /sn:0 /w:[ 0 ]
  //: input g10 (clk) @(739,507) /sn:0 /R:1 /w:[ 0 ]
  //: input g6 (Data) @(563,404) /sn:0 /w:[ 0 ]
  //: joint g7 (Reg2) @(454, 328) /w:[ 2 -1 1 4 ]
  //: output g9 (Data2) @(882,395) /sn:0 /w:[ 0 ]
  //: input g12 (clr) @(685,170) /sn:0 /w:[ 0 ]
  mux g5 (.I0(Reg2), .I1(RegMux), .S(RegDst), .Z(w12));   //: @(488,364) /sn:0 /R:1 /w:[ 5 1 1 0 ] /ss:0 /do:1
  //: input g11 (RegWrite) @(671,506) /sn:0 /R:1 /w:[ 0 ]
  //: input g14 (ESignExt) @(602,614) /sn:0 /w:[ 0 ]
  BRegs32x32 g0 (.clr(clr), .WriteData(Data), .Write(w12), .Read2(Reg2), .Read1(Reg1), .RegWrite(RegWrite), .clk(clk), .Data2(Data2), .Data1(Data1));   //: @(631, 256) /sz:(147, 182) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Li2>3 Li3>1 Bi0>1 Bi1>1 Ro0<1 Ro1<1 ]
  //: output g15 (SSignExt) @(822,613) /sn:0 /w:[ 1 ]
  SignExtend g13 (.E(ESignExt), .S(SSignExt));   //: @(658, 571) /sz:(93, 85) /sn:0 /p:[ Li0>1 Ro0<0 ]

endmodule

module SignExtend(S, E);
//: interface  /sz:(93, 85) /bd:[ Li0>E[15:0](43/85) Li1>E[15:0](43/85) Ro0<S[31:0](42/85) Ro1<S[31:0](42/85) ]
input [15:0] E;    //: /sn:0 {0}(225,137)(571,137)(571,155){1}
//: {2}(571,156)(571,165){3}
//: {4}(571,166)(571,175){5}
//: {6}(571,176)(571,185){7}
//: {8}(571,186)(571,195){9}
//: {10}(571,196)(571,205){11}
//: {12}(571,206)(571,215){13}
//: {14}(571,216)(571,225){15}
//: {16}(571,226)(571,235){17}
//: {18}(571,236)(571,245){19}
//: {20}(571,246)(571,255){21}
//: {22}(571,256)(571,265){23}
//: {24}(571,266)(571,275){25}
//: {26}(571,276)(571,285){27}
//: {28}(571,286)(571,295){29}
//: {30}(571,296)(571,305){31}
//: {32}(571,306)(571,315){33}
//: {34}(571,316)(571,325){35}
//: {36}(571,326)(571,335){37}
//: {38}(571,336)(571,345){39}
//: {40}(571,346)(571,355){41}
//: {42}(571,356)(571,365){43}
//: {44}(571,366)(571,375){45}
//: {46}(571,376)(571,385){47}
//: {48}(571,386)(571,395){49}
//: {50}(571,396)(571,405){51}
//: {52}(571,406)(571,415){53}
//: {54}(571,416)(571,425){55}
//: {56}(571,426)(571,435){57}
//: {58}(571,436)(571,445){59}
//: {60}(571,446)(571,455){61}
//: {62}(571,456)(571,465){63}
//: {64}(571,466)(571,501){65}
output [31:0] S;    //: /sn:0 {0}(881,311)(715,311){1}
wire w6;    //: /sn:0 {0}(709,396)(575,396){1}
wire w13;    //: /sn:0 {0}(709,326)(575,326){1}
wire w16;    //: /sn:0 {0}(709,296)(575,296){1}
wire w7;    //: /sn:0 {0}(709,386)(575,386){1}
wire w4;    //: /sn:0 {0}(709,416)(575,416){1}
wire w25;    //: /sn:0 {0}(709,206)(575,206){1}
wire w0;    //: /sn:0 {0}(709,446)(575,446){1}
wire w3;    //: /sn:0 {0}(709,426)(575,426){1}
wire w22;    //: /sn:0 {0}(709,236)(575,236){1}
wire w20;    //: /sn:0 {0}(709,256)(575,256){1}
wire w29;    //: /sn:0 {0}(709,166)(575,166){1}
wire w30;    //: /sn:0 {0}(709,156)(575,156){1}
wire w12;    //: /sn:0 {0}(709,336)(575,336){1}
wire w18;    //: /sn:0 {0}(709,276)(575,276){1}
wire w19;    //: /sn:0 {0}(709,266)(575,266){1}
wire w10;    //: /sn:0 {0}(709,356)(575,356){1}
wire w23;    //: /sn:0 {0}(709,226)(575,226){1}
wire w21;    //: /sn:0 {0}(709,246)(575,246){1}
wire w24;    //: /sn:0 {0}(709,216)(575,216){1}
wire w1;    //: /sn:0 {0}(709,436)(575,436){1}
wire w32;    //: /sn:0 {0}(575,456)(709,456){1}
wire w8;    //: /sn:0 {0}(709,376)(575,376){1}
wire w17;    //: /sn:0 {0}(709,286)(575,286){1}
wire w27;    //: /sn:0 {0}(709,186)(575,186){1}
wire w28;    //: /sn:0 {0}(709,176)(575,176){1}
wire w14;    //: /sn:0 {0}(709,316)(575,316){1}
wire w2;    //: /sn:0 {0}(575,466)(709,466){1}
wire w11;    //: /sn:0 {0}(709,346)(575,346){1}
wire w15;    //: /sn:0 {0}(709,306)(575,306){1}
wire w5;    //: /sn:0 {0}(709,406)(575,406){1}
wire w9;    //: /sn:0 {0}(709,366)(575,366){1}
wire w26;    //: /sn:0 {0}(709,196)(575,196){1}
//: enddecls

  tran g4(.Z(w32), .I(E[1]));   //: @(569,456) /sn:0 /R:2 /w:[ 0 62 61 ] /ss:1
  tran g8(.Z(w4), .I(E[5]));   //: @(569,416) /sn:0 /R:2 /w:[ 1 54 53 ] /ss:1
  concat g3 (.I0(w2), .I1(w32), .I2(w0), .I3(w1), .I4(w3), .I5(w4), .I6(w5), .I7(w6), .I8(w7), .I9(w8), .I10(w9), .I11(w10), .I12(w11), .I13(w12), .I14(w13), .I15(w14), .I16(w15), .I17(w16), .I18(w17), .I19(w18), .I20(w19), .I21(w20), .I22(w21), .I23(w22), .I24(w23), .I25(w24), .I26(w25), .I27(w26), .I28(w27), .I29(w28), .I30(w29), .I31(w30), .Z(S));   //: @(714,311) /sn:0 /w:[ 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0
  tran g16(.Z(w12), .I(E[13]));   //: @(569,336) /sn:0 /R:2 /w:[ 1 38 37 ] /ss:1
  tran g17(.Z(w13), .I(E[14]));   //: @(569,326) /sn:0 /R:2 /w:[ 1 36 35 ] /ss:1
  tran g26(.Z(w22), .I(E[15]));   //: @(569,236) /sn:0 /R:2 /w:[ 1 18 17 ] /ss:1
  tran g2(.Z(w2), .I(E[0]));   //: @(569,466) /sn:0 /R:2 /w:[ 0 64 63 ] /ss:1
  tran g23(.Z(w19), .I(E[15]));   //: @(569,266) /sn:0 /R:2 /w:[ 1 24 23 ] /ss:1
  tran g30(.Z(w26), .I(E[15]));   //: @(569,196) /sn:0 /R:2 /w:[ 1 10 9 ] /ss:1
  //: output g1 (S) @(878,311) /sn:0 /w:[ 0 ]
  tran g24(.Z(w20), .I(E[15]));   //: @(569,256) /sn:0 /R:2 /w:[ 1 22 21 ] /ss:1
  tran g29(.Z(w25), .I(E[15]));   //: @(569,206) /sn:0 /R:2 /w:[ 1 12 11 ] /ss:1
  tran g18(.Z(w14), .I(E[15]));   //: @(569,316) /sn:0 /R:2 /w:[ 1 34 33 ] /ss:1
  tran g10(.Z(w6), .I(E[7]));   //: @(569,396) /sn:0 /R:2 /w:[ 1 50 49 ] /ss:1
  tran g25(.Z(w21), .I(E[15]));   //: @(569,246) /sn:0 /R:2 /w:[ 1 20 19 ] /ss:1
  tran g6(.Z(w1), .I(E[3]));   //: @(569,436) /sn:0 /R:2 /w:[ 1 58 57 ] /ss:1
  tran g7(.Z(w3), .I(E[4]));   //: @(569,426) /sn:0 /R:2 /w:[ 1 56 55 ] /ss:1
  tran g9(.Z(w5), .I(E[6]));   //: @(569,406) /sn:0 /R:2 /w:[ 1 52 51 ] /ss:1
  tran g22(.Z(w18), .I(E[15]));   //: @(569,276) /sn:0 /R:2 /w:[ 1 26 25 ] /ss:1
  tran g31(.Z(w27), .I(E[15]));   //: @(569,186) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  tran g33(.Z(w29), .I(E[15]));   //: @(569,166) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  tran g12(.Z(w8), .I(E[9]));   //: @(569,376) /sn:0 /R:2 /w:[ 1 46 45 ] /ss:1
  tran g28(.Z(w24), .I(E[15]));   //: @(569,216) /sn:0 /R:2 /w:[ 1 14 13 ] /ss:1
  tran g34(.Z(w30), .I(E[15]));   //: @(569,156) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  tran g5(.Z(w0), .I(E[2]));   //: @(569,446) /sn:0 /R:2 /w:[ 1 60 59 ] /ss:1
  tran g11(.Z(w7), .I(E[8]));   //: @(569,386) /sn:0 /R:2 /w:[ 1 48 47 ] /ss:1
  tran g14(.Z(w10), .I(E[11]));   //: @(569,356) /sn:0 /R:2 /w:[ 1 42 41 ] /ss:1
  tran g19(.Z(w15), .I(E[15]));   //: @(569,306) /sn:0 /R:2 /w:[ 1 32 31 ] /ss:1
  tran g21(.Z(w17), .I(E[15]));   //: @(569,286) /sn:0 /R:2 /w:[ 1 28 27 ] /ss:1
  tran g20(.Z(w16), .I(E[15]));   //: @(569,296) /sn:0 /R:2 /w:[ 1 30 29 ] /ss:1
  tran g32(.Z(w28), .I(E[15]));   //: @(569,176) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  //: input g0 (E) @(223,137) /sn:0 /w:[ 0 ]
  tran g15(.Z(w11), .I(E[12]));   //: @(569,346) /sn:0 /R:2 /w:[ 1 40 39 ] /ss:1
  tran g27(.Z(w23), .I(E[15]));   //: @(569,226) /sn:0 /R:2 /w:[ 1 16 15 ] /ss:1
  tran g13(.Z(w9), .I(E[10]));   //: @(569,366) /sn:0 /R:2 /w:[ 1 44 43 ] /ss:1

endmodule

module FormatoI(RegDst, Zero, Inst, MemWrite, RegWrite, MemtoReg, clr, ALUSrc, clk, MemRead, ALUOp);
//: interface  /sz:(40, 40) /bd:[ ]
input Zero;    //: /sn:0 {0}(1059,290)(1009,290){1}
input MemWrite;    //: /sn:0 {0}(1204,224)(1204,259){1}
input ALUSrc;    //: /sn:0 {0}(719,449)(719,396){1}
input [31:0] Inst;    //: /sn:0 {0}(236,173)(236,242){1}
//: {2}(236,243)(236,284){3}
//: {4}(236,285)(236,328){5}
//: {6}(236,329)(236,418){7}
//: {8}(236,419)(236,509){9}
input RegDst;    //: /sn:0 {0}(308,368)(359,368){1}
input clr;    //: /sn:0 {0}(491,186)(491,215){1}
input RegWrite;    //: /sn:0 {0}(476,520)(476,464){1}
input clk;    //: /sn:0 {0}(520,537)(520,510){1}
input [3:0] ALUOp;    //: /sn:0 {0}(855,197)(855,240){1}
input MemtoReg;    //: /sn:0 {0}(1387,479)(1387,437){1}
input MemRead;    //: /sn:0 {0}(1202,498)(1202,460){1}
wire w6;    //: /sn:0 {0}(520,494)(520,464){1}
wire [31:0] w7;    //: /sn:0 /dp:1 {0}(1371,404)(1314,404)(1314,356)(1264,356){1}
wire [4:0] w4;    //: /sn:0 {0}(359,293)(248,293)(248,285)(240,285){1}
wire [31:0] w0;    //: /sn:0 /dp:1 {0}(703,383)(655,383)(655,412)(605,412){1}
wire [4:0] w3;    //: /sn:0 {0}(359,333)(248,333)(248,329)(240,329){1}
wire [31:0] w18;    //: /sn:0 {0}(1134,426)(682,426)(682,365){1}
//: {2}(684,363)(703,363){3}
//: {4}(680,363)(653,363)(653,342)(605,342){5}
wire [31:0] w10;    //: /sn:0 {0}(1400,414)(1410,414)(1410,572)(422,572)(422,464){1}
wire [15:0] w1;    //: /sn:0 {0}(359,418)(248,418)(248,419)(240,419){1}
wire [31:0] w14;    //: /sn:0 {0}(732,373)(793,373)(793,342)(801,342){1}
wire [31:0] w11;    //: /sn:0 {0}(605,279)(801,279){1}
wire [31:0] w15;    //: /sn:0 {0}(1009,330)(1064,330){1}
//: {2}(1068,330)(1134,330){3}
//: {4}(1066,332)(1066,528)(1315,528)(1315,424)(1371,424){5}
wire [4:0] w5;    //: /sn:0 {0}(359,247)(248,247)(248,243)(240,243){1}
//: enddecls

  //: input g8 (RegDst) @(306,368) /sn:0 /w:[ 0 ]
  tran g4(.Z(w1), .I(Inst[15:0]));   //: @(234,419) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  //: input g16 (Zero) @(1061,290) /sn:0 /R:2 /w:[ 0 ]
  //: input g3 (Inst) @(236,171) /sn:0 /R:3 /w:[ 0 ]
  //: input g17 (MemWrite) @(1204,222) /sn:0 /R:3 /w:[ 0 ]
  MEM g2 (.MemWrite(MemWrite), .Address(w15), .WriteData(w18), .MemRead(MemRead), .ReadData(w7));   //: @(1135, 260) /sz:(128, 199) /sn:0 /p:[ Ti0>1 Li0>3 Li1>0 Bi0>1 Ro0<1 ]
  ALU g1 (.ALUOp(ALUOp), .A(w11), .B(w14), .Zero(Zero), .ALURes(w15));   //: @(802, 241) /sz:(206, 161) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  //: joint g18 (w18) @(682, 363) /w:[ 2 -1 4 1 ]
  not g10 (.I(clk), .Z(w6));   //: @(520,504) /sn:0 /R:1 /w:[ 1 0 ]
  tran g6(.Z(w4), .I(Inst[4:0]));   //: @(234,285) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  //: input g9 (RegWrite) @(476,522) /sn:0 /R:1 /w:[ 0 ]
  tran g7(.Z(w5), .I(Inst[4:0]));   //: @(234,243) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  //: input g22 (MemtoReg) @(1387,481) /sn:0 /R:1 /w:[ 0 ]
  //: input g12 (clr) @(491,184) /sn:0 /R:3 /w:[ 0 ]
  //: input g14 (ALUSrc) @(719,451) /sn:0 /R:1 /w:[ 0 ]
  //: input g11 (clk) @(520,539) /sn:0 /R:1 /w:[ 0 ]
  tran g5(.Z(w3), .I(Inst[4:0]));   //: @(234,329) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  //: joint g21 (w15) @(1066, 330) /w:[ 2 -1 1 4 ]
  //: input g19 (MemRead) @(1202,500) /sn:0 /R:1 /w:[ 0 ]
  mux g20 (.I0(w15), .I1(w7), .S(MemtoReg), .Z(w10));   //: @(1387,414) /sn:0 /R:1 /w:[ 5 0 1 0 ] /ss:0 /do:0
  //: input g15 (ALUOp) @(855,195) /sn:0 /R:3 /w:[ 0 ]
  READ g0 (.clr(clr), .Reg1(w5), .Reg2(w4), .RegMux(w3), .RegDst(RegDst), .ESignExt(w1), .Data(w10), .clk(w6), .RegWrite(RegWrite), .Data1(w11), .Data2(w18), .SSignExt(w0));   //: @(360, 216) /sz:(244, 247) /sn:0 /p:[ Ti0>1 Li0>0 Li1>0 Li2>0 Li3>1 Li4>0 Bi0>1 Bi1>1 Bi2>1 Ro0<0 Ro1<5 Ro2<1 ]
  mux g13 (.I0(w0), .I1(w18), .S(ALUSrc), .Z(w14));   //: @(719,373) /sn:0 /R:1 /w:[ 0 3 1 0 ] /ss:0 /do:0

endmodule

module ALU(ALURes, Zero, ALUOp, B, A);
//: interface  /sz:(206, 161) /bd:[ Ti0>ALUOp[3:0](53/206) Ti1>ALUOp[3:0](53/206) Li0>A[31:0](38/161) Li1>B[31:0](101/161) Li2>B[31:0](101/161) Li3>A[31:0](38/161) Ro0<Zero(49/161) Ro1<ALURes[31:0](109/161) Ro2<ALURes[31:0](89/161) Ro3<Zero(49/161) ]
input [31:0] B;    //: /sn:0 {0}(463,286)(453,286)(453,296)(397,296)(397,251){1}
//: {2}(399,249)(455,249)(455,230)(465,230){3}
//: {4}(395,249)(346,249){5}
//: {6}(342,249)(288,249){7}
//: {8}(284,249)(226,249){9}
//: {10}(286,251)(286,462)(354,462){11}
//: {12}(344,251)(344,370)(459,370){13}
output Zero;    //: /sn:0 /dp:1 {0}(820,634)(868,634){1}
input [31:0] A;    //: /sn:0 {0}(228,202)(311,202){1}
//: {2}(315,202)(370,202){3}
//: {4}(374,202)(409,202){5}
//: {6}(413,202)(456,202)(456,225)(465,225){7}
//: {8}(411,204)(411,270)(453,270)(453,281)(463,281){9}
//: {10}(372,204)(372,338)(459,338){11}
//: {12}(313,204)(313,430)(459,430){13}
supply0 w0;    //: /sn:0 {0}(493,315)(473,315)(473,330){1}
supply1 w1;    //: /sn:0 {0}(499,401)(473,401)(473,422){1}
input [3:0] ALUOp;    //: /sn:0 /dp:3 {0}(633,620)(633,596){1}
//: {2}(633,595)(633,574)(626,574){3}
output [31:0] ALURes;    //: /sn:0 {0}(746,609)(746,669)(770,669){1}
//: {2}(774,669)(792,669)(792,700){3}
//: {4}(772,667)(772,634)(799,634){5}
wire [31:0] w16;    //: /sn:0 {0}(370,462)(459,462){1}
wire [31:0] w7;    //: /sn:0 {0}(943,512)(943,560)(766,560)(766,580){1}
wire [31:0] w4;    //: /sn:0 {0}(484,283)(736,283)(736,580){1}
wire [2:0] w3;    //: /sn:0 /dp:1 {0}(637,596)(723,596){1}
wire [31:0] w12;    //: /sn:0 {0}(488,446)(754,446){1}
//: {2}(758,446)(943,446)(943,491){3}
//: {4}(756,448)(756,580){5}
wire [31:0] w10;    //: /sn:0 {0}(488,354)(746,354)(746,580){1}
wire w14;    //: /sn:0 {0}(473,470)(473,480){1}
wire [31:0] w2;    //: /sn:0 {0}(486,228)(726,228)(726,580){1}
wire [4:0] w15;    //: /sn:0 /dp:1 {0}(859,482)(859,501)(906,501){1}
wire Zero0;    //: /sn:0 {0}(473,378)(473,385){1}
//: enddecls

  //: joint g8 (B) @(397, 249) /w:[ 2 -1 4 1 ]
  //: output g4 (ALURes) @(792,697) /sn:0 /R:3 /w:[ 3 ]
  //: joint g16 (A) @(313, 202) /w:[ 2 -1 1 12 ]
  //: output g3 (Zero) @(865,634) /sn:0 /w:[ 1 ]
  //: supply0 g17 (w0) @(499,315) /sn:0 /R:1 /w:[ 0 ]
  //: input g2 (ALUOp) @(624,574) /sn:0 /w:[ 3 ]
  //: joint g23 (ALURes) @(772, 669) /w:[ 2 4 1 -1 ]
  //: input g1 (B) @(224,249) /sn:0 /w:[ 9 ]
  tran g24(.Z(w3), .I(ALUOp[2:0]));   //: @(631,596) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  //: supply1 g18 (w1) @(499,412) /sn:0 /R:3 /w:[ 0 ]
  add g10 (.A(B), .B(A), .S(w10), .CI(w0), .CO(Zero0));   //: @(475,354) /sn:0 /R:1 /w:[ 13 11 0 1 0 ]
  or g6 (.I0(A), .I1(B), .Z(w4));   //: @(474,283) /sn:0 /w:[ 9 0 0 ]
  mux g9 (.I0(w2), .I1(w4), .I2(w10), .I3(w12), .I4(w7), .S(w3), .Z(ALURes));   //: @(746,596) /sn:0 /w:[ 1 1 1 5 1 1 0 ] /ss:0 /do:0
  //: joint g7 (A) @(411, 202) /w:[ 6 -1 5 8 ]
  //: dip g22 (w15) @(859,472) /sn:0 /w:[ 0 ] /st:31
  //: joint g12 (B) @(344, 249) /w:[ 5 -1 6 12 ]
  not g14 (.I(B), .Z(w16));   //: @(360,462) /sn:0 /w:[ 11 0 ]
  //: joint g11 (A) @(372, 202) /w:[ 4 -1 3 10 ]
  and g5 (.I0(A), .I1(B), .Z(w2));   //: @(476,228) /sn:0 /w:[ 7 3 0 ]
  nor g19 (.I0(ALURes), .Z(Zero));   //: @(810,634) /sn:0 /w:[ 5 0 ]
  rshift g21 (.I(w12), .Z(w7), .S(w15));   //: @(943,501) /sn:0 /w:[ 3 0 1 ]
  //: joint g20 (w12) @(756, 446) /w:[ 2 -1 1 4 ]
  //: joint g15 (B) @(286, 249) /w:[ 7 -1 8 10 ]
  //: input g0 (A) @(226,202) /sn:0 /w:[ 0 ]
  add g13 (.A(w16), .B(A), .S(w12), .CI(w1), .CO(w14));   //: @(475,446) /sn:0 /R:1 /w:[ 1 13 0 1 0 ]

endmodule

module BRegs32x32(Read2, Write, Read1, Data2, Data1, clr, clk, RegWrite, WriteData);
//: interface  /sz:(147, 182) /bd:[ Ti0>clr(66/147) Ti1>clr(66/147) Li0>Read1[4:0](32/182) Li1>Read2[4:0](72/182) Li2>Write[4:0](108/182) Li3>WriteData[31:0](148/182) Li4>WriteData[31:0](148/182) Li5>Write[4:0](108/182) Li6>Read2[4:0](72/182) Li7>Read1[4:0](32/182) Bi0>clk(108/147) Bi1>RegWrite(40/147) Bi2>RegWrite(40/147) Bi3>clk(108/147) Ro0<Data1[31:0](47/182) Ro1<Data2[31:0](139/182) Ro2<Data2[31:0](139/182) Ro3<Data1[31:0](47/182) ]
output [31:0] Data2;    //: /sn:0 {0}(668,485)(668,472)(669,472)(669,445){1}
input [4:0] Write;    //: /sn:0 {0}(-238,-38)(-138,-38)(-138,-37)(-66,-37){1}
//: {2}(-65,-37)(-28,-37){3}
//: {4}(-27,-37)(-16,-37){5}
input [31:0] WriteData;    //: /sn:0 {0}(669,157)(669,75)(481,75){1}
//: {2}(477,75)(292,75){3}
//: {4}(288,75)(89,75){5}
//: {6}(85,75)(-104,75)(-104,73)(-237,73){7}
//: {8}(87,77)(87,157){9}
//: {10}(290,77)(290,107)(291,107)(291,152){11}
//: {12}(479,77)(479,157){13}
supply1 w21;    //: /sn:0 {0}(82,3)(57,3)(57,-11){1}
output [31:0] Data1;    //: /sn:0 {0}(59,382)(59,465){1}
input RegWrite;    //: /sn:0 {0}(-237,263)(-71,263){1}
//: {2}(-67,263)(171,263){3}
//: {4}(175,263)(370,263){5}
//: {6}(374,263)(552,263)(552,219)(556,219){7}
//: {8}(372,261)(372,219)(383,219){9}
//: {10}(173,261)(173,214)(183,214){11}
//: {12}(-69,261)(-69,219)(-38,219){13}
input clr;    //: /sn:0 {0}(721,193)(731,193)(731,-83)(543,-83){1}
//: {2}(539,-83)(355,-83){3}
//: {4}(351,-83)(150,-83){5}
//: {6}(146,-83)(-44,-83)(-44,-92)(-235,-92){7}
//: {8}(148,-81)(148,193)(139,193){9}
//: {10}(353,-81)(353,188)(343,188){11}
//: {12}(541,-81)(541,193)(531,193){13}
input clk;    //: /sn:0 {0}(556,214)(542,214)(542,285)(364,285){1}
//: {2}(362,283)(362,214)(383,214){3}
//: {4}(360,285)(167,285){5}
//: {6}(165,283)(165,209)(183,209){7}
//: {8}(163,285)(-56,285){9}
//: {10}(-58,283)(-58,214)(-38,214){11}
//: {12}(-60,285)(-237,285){13}
input [4:0] Read1;    //: {0}(-237,96)(-208,96)(-208,95)(-124,95){1}
//: {2}(-123,95)(-96,95){3}
//: {4}(-95,95)(-78,95){5}
input [4:0] Read2;    //: {0}(-237,145)(-141,145){1}
//: {2}(-140,145)(-123,145)(-123,144)(-94,144){3}
//: {4}(-93,144)(-79,144){5}
wire w16;    //: /sn:0 {0}(39,205)(-50,205)(-50,39)(88,39)(88,19){1}
wire [1:0] w6;    //: /sn:0 {0}(36,369)(-123,369)(-123,99){1}
wire w4;    //: /sn:0 {0}(112,19)(112,46)(370,46)(370,205)(431,205){1}
wire w22;    //: /sn:0 {0}(404,217)(431,217){1}
wire [31:0] w0;    //: /sn:0 {0}(651,416)(651,398)(105,398)(105,228){1}
wire [31:0] R2;    //: {0}(65,353)(65,319)(469,319)(469,228){1}
wire [31:0] w3;    //: /sn:0 {0}(77,353)(77,334)(659,334)(659,228){1}
wire w20;    //: /sn:0 {0}(124,19)(124,29)(556,29)(556,205)(621,205){1}
wire [2:0] w18;    //: /sn:0 {0}(431,180)(402,180)(402,125){1}
//: {2}(404,123)(589,123)(589,180)(621,180){3}
//: {4}(400,123)(279,123)(279,122)(212,122){5}
//: {6}(208,122)(8,122){7}
//: {8}(4,122)(-93,122)(-93,139){9}
//: {10}(6,124)(6,180)(39,180){11}
//: {12}(210,124)(210,175)(243,175){13}
wire [2:0] w19;    //: /sn:0 {0}(431,169)(419,169)(419,109){1}
//: {2}(421,107)(606,107)(606,169)(621,169){3}
//: {4}(417,107)(297,107)(297,106)(231,106){5}
//: {6}(227,106)(25,106){7}
//: {8}(21,106)(-95,106)(-95,99){9}
//: {10}(23,108)(23,169)(39,169){11}
//: {12}(229,108)(229,164)(243,164){13}
wire [1:0] w10;    //: /sn:0 {0}(-140,149)(-140,432)(646,432){1}
wire w23;    //: /sn:0 {0}(577,217)(621,217){1}
wire [2:0] w24;    //: /sn:0 {0}(431,193)(381,193)(381,141){1}
//: {2}(383,139)(568,139)(568,193)(621,193){3}
//: {4}(379,139)(260,139)(260,138)(195,138){5}
//: {6}(191,138)(-13,138){7}
//: {8}(-17,138)(-65,138)(-65,-33){9}
//: {10}(-15,140)(-15,193)(39,193){11}
//: {12}(193,140)(193,188)(243,188){13}
wire w1;    //: /sn:0 {0}(-17,217)(39,217){1}
wire w31;    //: /sn:0 {0}(243,200)(178,200)(178,60)(100,60)(100,19){1}
wire [31:0] R3;    //: {0}(687,228)(687,416){1}
wire [31:0] R1;    //: {0}(281,223)(281,308)(53,308)(53,353){1}
wire w2;    //: /sn:0 {0}(243,212)(204,212){1}
wire [1:0] w11;    //: /sn:0 {0}(-27,-33)(-27,-23)(106,-23)(106,-10){1}
wire [31:0] R0;    //: {0}(77,228)(77,299)(41,299)(41,353){1}
wire [31:0] w5;    //: /sn:0 {0}(675,416)(675,372)(497,372)(497,228){1}
wire [31:0] w9;    //: /sn:0 {0}(663,416)(663,387)(309,387)(309,223){1}
//: enddecls

  //: joint g44 (clr) @(353, -83) /w:[ 3 -1 4 10 ]
  //: input g4 (Read2) @(-239,145) /sn:0 /w:[ 0 ]
  //: joint g8 (w18) @(6, 122) /w:[ 7 -1 8 10 ]
  //: joint g47 (clr) @(541, -83) /w:[ 1 -1 2 12 ]
  //: joint g16 (clk) @(165, 285) /w:[ 5 6 8 -1 ]
  //: input g3 (Write) @(-240,-38) /sn:0 /w:[ 0 ]
  //: joint g26 (w19) @(229, 106) /w:[ 5 -1 6 12 ]
  //: input g17 (Read1) @(-239,96) /sn:0 /w:[ 0 ]
  //: output g2 (Data2) @(668,482) /sn:0 /R:3 /w:[ 0 ]
  tran g30(.Z(w10), .I(Read2[4:3]));   //: @(-140,143) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g23(.Z(w24), .I(Write[2:0]));   //: @(-65,-39) /sn:0 /R:1 /w:[ 9 1 2 ] /ss:1
  Regs8x32 g24 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w31), .clk(w2), .clr(clr), .AOUT(R1), .BOUT(w9));   //: @(244, 153) /sz:(98, 69) /sn:0 /p:[ Ti0>11 Li0>13 Li1>13 Li2>13 Li3>0 Li4>0 Ri0>11 Bo0<0 Bo1<1 ]
  //: joint g39 (RegWrite) @(372, 263) /w:[ 6 8 5 -1 ]
  //: output g1 (Data1) @(59,462) /sn:0 /R:3 /w:[ 1 ]
  Regs8x32 g29 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w4), .clk(w22), .clr(clr), .AOUT(R2), .BOUT(w5));   //: @(432, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>13 Li0>0 Li1>0 Li2>0 Li3>1 Li4>1 Ri0>13 Bo0<1 Bo1<1 ]
  //: comment g51 /dolink:0 /link:"" @(395,229) /sn:0
  //: /line:"Regs 16-23"
  //: /end
  tran g18(.Z(w19), .I(Read1[2:0]));   //: @(-95,93) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:1
  //: joint g25 (w18) @(210, 122) /w:[ 5 -1 6 12 ]
  //: supply1 g10 (w21) @(68,-11) /sn:0 /w:[ 1 ]
  //: comment g49 /dolink:0 /link:"" @(210,225) /sn:0
  //: /line:"Regs 8-15"
  //: /end
  Regs8x32 g6 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w16), .clk(w1), .clr(clr), .AOUT(R0), .BOUT(w0));   //: @(40, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>9 Li0>11 Li1>11 Li2>11 Li3>0 Li4>1 Ri0>9 Bo0<0 Bo1<1 ]
  //: comment g50 /dolink:0 /link:"" @(585,229) /sn:0
  //: /line:"Regs 24-31"
  //: /end
  and g35 (.I0(clk), .I1(RegWrite), .Z(w22));   //: @(394,217) /sn:0 /delay:" 1" /w:[ 3 9 0 ]
  demux g9 (.I(w11), .E(w21), .Z0(w16), .Z1(w31), .Z2(w4), .Z3(w20));   //: @(106,3) /sn:0 /w:[ 1 0 1 1 0 0 ]
  //: joint g7 (w19) @(23, 106) /w:[ 7 -1 8 10 ]
  tran g22(.Z(w18), .I(Read2[2:0]));   //: @(-93,142) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:0
  tran g31(.Z(w6), .I(Read1[4:3]));   //: @(-123,93) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  and g33 (.I0(clk), .I1(RegWrite), .Z(w1));   //: @(-27,217) /sn:0 /delay:" 1" /w:[ 11 13 0 ]
  //: joint g45 (WriteData) @(479, 75) /w:[ 1 -1 2 12 ]
  //: joint g41 (w19) @(419, 107) /w:[ 2 -1 4 1 ]
  and g36 (.I0(clk), .I1(RegWrite), .Z(w23));   //: @(567,217) /sn:0 /delay:" 1" /w:[ 0 7 0 ]
  //: joint g40 (w18) @(402, 123) /w:[ 2 -1 4 1 ]
  //: input g42 (clr) @(-237,-92) /sn:0 /w:[ 7 ]
  //: input g12 (clk) @(-239,285) /sn:0 /w:[ 13 ]
  Regs8x32 g46 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w20), .clk(w23), .clr(clr), .AOUT(w3), .BOUT(R3));   //: @(622, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>0 Li0>3 Li1>3 Li2>3 Li3>1 Li4>1 Ri0>0 Bo0<1 Bo1<0 ]
  //: joint g28 (w24) @(381, 139) /w:[ 2 -1 4 1 ]
  and g34 (.I0(clk), .I1(RegWrite), .Z(w2));   //: @(194,212) /sn:0 /delay:" 1" /w:[ 7 11 1 ]
  tran g5(.Z(w11), .I(Write[4:3]));   //: @(-27,-39) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  mux g14 (.I0(R0), .I1(R1), .I2(R2), .I3(w3), .S(w6), .Z(Data1));   //: @(59,369) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  //: joint g11 (w24) @(-15, 138) /w:[ 7 -1 8 10 ]
  //: joint g21 (w24) @(193, 138) /w:[ 5 -1 6 12 ]
  //: joint g19 (clk) @(-58, 285) /w:[ 9 10 12 -1 ]
  //: joint g20 (WriteData) @(87, 75) /w:[ 5 -1 6 8 ]
  //: input g32 (RegWrite) @(-239,263) /sn:0 /w:[ 0 ]
  //: input g0 (WriteData) @(-239,73) /sn:0 /w:[ 7 ]
  //: joint g43 (clr) @(148, -83) /w:[ 5 -1 6 8 ]
  //: joint g15 (clk) @(362, 285) /w:[ 1 2 4 -1 ]
  //: joint g38 (RegWrite) @(173, 263) /w:[ 4 10 3 -1 ]
  //: comment g48 /dolink:0 /link:"" @(11,228) /sn:0
  //: /line:"Regs 0-7"
  //: /end
  //: joint g27 (WriteData) @(290, 75) /w:[ 3 -1 4 10 ]
  //: joint g37 (RegWrite) @(-69, 263) /w:[ 2 12 1 -1 ]
  mux g13 (.I0(w0), .I1(w9), .I2(w5), .I3(R3), .S(w10), .Z(Data2));   //: @(669,432) /sn:0 /w:[ 0 0 0 1 1 1 ] /ss:0 /do:0

endmodule

module Regs8x32(SB, SA, BOUT, AOUT, clr, clk, RegWr, SD, DIN);
//: interface  /sz:(98, 69) /bd:[ Ti0>DIN[31:0](47/98) Ti1>DIN[31:0](47/98) Ti2>DIN[31:0](47/98) Ti3>DIN[31:0](47/98) Li0>SD[2:0](35/69) Li1>SA[2:0](11/69) Li2>SB[2:0](22/69) Li3>RegWr(47/69) Li4>clk(59/69) Li5>SD[2:0](35/69) Li6>SA[2:0](11/69) Li7>SB[2:0](22/69) Li8>RegWr(47/69) Li9>clk(59/69) Li10>clk(59/69) Li11>RegWr(47/69) Li12>SB[2:0](22/69) Li13>SA[2:0](11/69) Li14>SD[2:0](35/69) Li15>clk(59/69) Li16>RegWr(47/69) Li17>SB[2:0](22/69) Li18>SA[2:0](11/69) Li19>SD[2:0](35/69) Ri0>clr(35/69) Ri1>clr(35/69) Ri2>clr(35/69) Ri3>clr(35/69) Bo0<AOUT[31:0](37/98) Bo1<BOUT[31:0](65/98) Bo2<AOUT[31:0](37/98) Bo3<BOUT[31:0](65/98) Bo4<BOUT[31:0](65/98) Bo5<AOUT[31:0](37/98) Bo6<BOUT[31:0](65/98) Bo7<AOUT[31:0](37/98) ]
input [31:0] DIN;    //: /sn:0 {0}(531,269)(531,318){1}
//: {2}(533,320)(627,320){3}
//: {4}(631,320)(715,320){5}
//: {6}(719,320)(807,320)(807,429){7}
//: {8}(717,322)(717,352){9}
//: {10}(629,322)(629,433){11}
//: {12}(529,320)(435,320){13}
//: {14}(431,320)(342,320){15}
//: {16}(338,320)(264,320){17}
//: {18}(260,320)(181,320)(181,352){19}
//: {20}(262,322)(262,439){21}
//: {22}(340,322)(340,351){23}
//: {24}(433,322)(433,436){25}
//: {26}(531,322)(531,348){27}
output [31:0] BOUT;    //: /sn:0 {0}(516,697)(516,672){1}
input [2:0] SD;    //: /sn:0 {0}(782,138)(852,138)(852,156){1}
input [2:0] SB;    //: /sn:0 {0}(466,659)(493,659){1}
supply1 w21;    //: /sn:0 {0}(828,169)(801,169)(801,153){1}
input RegWr;    //: /sn:0 {0}(48,363)(68,363)(68,378)(82,378){1}
input clr;    //: /sn:0 /dp:1 {0}(959,337)(1032,337){1}
input [2:0] SA;    //: /sn:0 {0}(256,657)(231,657){1}
input clk;    //: /sn:0 {0}(82,383)(68,383)(68,398)(55,398){1}
output [31:0] AOUT;    //: /sn:0 {0}(279,670)(279,702){1}
wire [31:0] w16;    //: /sn:0 {0}(531,369)(531,574)(520,574){1}
//: {2}(516,574)(282,574)(282,641){3}
//: {4}(518,576)(518,587)(519,587)(519,643){5}
wire w7;    //: /sn:0 {0}(472,451)(513,451)(513,405)(848,405)(848,185){1}
wire [31:0] R5;    //: {0}(288,641)(288,586)(525,586){1}
//: {2}(529,586)(629,586)(629,454){3}
//: {4}(527,588)(527,617)(525,617)(525,643){5}
wire w4;    //: /sn:0 {0}(943,337)(906,337){1}
//: {2}(902,337)(767,337){3}
//: {4}(763,337)(588,337){5}
//: {6}(584,337)(390,337){7}
//: {8}(386,337)(231,337)(231,357)(220,357){9}
//: {10}(388,339)(388,356)(379,356){11}
//: {12}(586,339)(586,353)(570,353){13}
//: {14}(765,339)(765,357)(756,357){15}
//: {16}(904,339)(904,417)(865,417){17}
//: {18}(861,417)(675,417){19}
//: {20}(671,417)(489,417){21}
//: {22}(485,417)(302,417)(302,444)(301,444){23}
//: {24}(487,419)(487,441)(472,441){25}
//: {26}(673,419)(673,438)(668,438){27}
//: {28}(863,419)(863,434)(846,434){29}
wire w3;    //: /sn:0 {0}(835,185)(835,397)(330,397)(330,454)(301,454){1}
wire w0;    //: /sn:0 {0}(770,439)(764,439)(764,481)(579,481){1}
//: {2}(577,479)(577,443)(592,443){3}
//: {4}(575,481)(390,481){5}
//: {6}(388,479)(388,446)(396,446){7}
//: {8}(386,481)(214,481){9}
//: {10}(212,479)(212,449)(225,449){11}
//: {12}(210,481)(125,481)(125,383){13}
//: {14}(127,381)(291,381){15}
//: {16}(295,381)(477,381){17}
//: {18}(481,381)(660,381)(660,362)(680,362){19}
//: {20}(479,379)(479,358)(494,358){21}
//: {22}(293,379)(293,361)(303,361){23}
//: {24}(125,379)(125,362)(144,362){25}
//: {26}(123,381)(103,381){27}
wire [31:0] R2;    //: {0}(262,641)(262,537){1}
//: {2}(264,535)(499,535)(499,643){3}
//: {4}(262,533)(262,460){5}
wire [31:0] R7;    //: {0}(807,450)(807,609)(541,609){1}
//: {2}(537,609)(302,609)(302,641){3}
//: {4}(539,611)(539,643){5}
wire w12;    //: /sn:0 {0}(756,367)(787,367)(787,258)(868,258)(868,185){1}
wire w10;    //: /sn:0 {0}(846,444)(875,444)(875,185){1}
wire [31:0] R4;    //: {0}(340,372)(340,545){1}
//: {2}(342,547)(505,547)(505,643){3}
//: {4}(338,547)(268,547)(268,641){5}
wire [31:0] R3;    //: {0}(512,643)(512,559)(435,559){1}
//: {2}(433,557)(433,457){3}
//: {4}(431,559)(275,559)(275,641){5}
wire w8;    //: /sn:0 {0}(220,367)(249,367)(249,213)(828,213)(828,185){1}
wire Z5;    //: /sn:0 {0}(861,185)(861,413)(700,413)(700,448)(668,448){1}
wire w14;    //: /sn:0 {0}(379,366)(414,366)(414,229)(841,229)(841,185){1}
wire [31:0] R0;    //: {0}(492,643)(492,523)(257,523){1}
//: {2}(253,523)(181,523)(181,373){3}
//: {4}(255,525)(255,641){5}
wire w15;    //: /sn:0 {0}(570,363)(608,363)(608,244)(855,244)(855,185){1}
wire [31:0] R10;    //: /sn:0 {0}(295,641)(295,600)(530,600){1}
//: {2}(534,600)(717,600)(717,373){3}
//: {4}(532,602)(532,643){5}
//: enddecls

  //: input g4 (SB) @(464,659) /sn:0 /w:[ 0 ]
  //: joint g8 (w16) @(518, 574) /w:[ 1 -1 2 4 ]
  //: joint g16 (R3) @(433, 559) /w:[ 1 2 4 -1 ]
  //: input g3 (SA) @(229,657) /sn:0 /w:[ 1 ]
  //: joint g26 (DIN) @(340, 320) /w:[ 15 -1 16 22 ]
  //: joint g17 (R4) @(340, 547) /w:[ 2 1 4 -1 ]
  //: output g2 (BOUT) @(516,694) /sn:0 /R:3 /w:[ 0 ]
  register R5 (.Q(R5), .D(DIN), .EN(Z5), .CLR(w4), .CK(!w0));   //: @(629,443) /w:[ 3 11 1 27 3 ]
  //: joint g30 (w0) @(212, 481) /w:[ 9 10 12 -1 ]
  //: joint g23 (w4) @(765, 337) /w:[ 3 -1 4 14 ]
  //: joint g24 (DIN) @(531, 320) /w:[ 2 1 12 26 ]
  //: joint g39 (DIN) @(262, 320) /w:[ 17 -1 18 20 ]
  //: output g1 (AOUT) @(279,699) /sn:0 /R:3 /w:[ 1 ]
  //: joint g29 (w0) @(388, 481) /w:[ 5 6 8 -1 ]
  register R2 (.Q(R4), .D(DIN), .EN(w14), .CLR(w4), .CK(!w0));   //: @(340,361) /w:[ 0 23 0 11 23 ]
  //: joint g18 (R2) @(262, 535) /w:[ 2 4 -1 1 ]
  register R7 (.Q(R7), .D(DIN), .EN(w10), .CLR(w4), .CK(!w0));   //: @(807,439) /w:[ 0 7 0 29 0 ]
  not g25 (.I(clr), .Z(w4));   //: @(953,337) /sn:0 /R:2 /w:[ 0 0 ]
  //: supply1 g10 (w21) @(812,153) /sn:0 /w:[ 1 ]
  register R6 (.Q(R10), .D(DIN), .EN(w12), .CLR(w4), .CK(!w0));   //: @(717,362) /w:[ 3 9 0 15 19 ]
  //: joint g6 (R7) @(539, 609) /w:[ 1 -1 2 4 ]
  and g35 (.I0(RegWr), .I1(clk), .Z(w0));   //: @(93,381) /sn:0 /delay:" 1" /w:[ 1 0 27 ]
  demux g9 (.I(SD), .E(w21), .Z0(!w8), .Z1(!w3), .Z2(!w14), .Z3(!w7), .Z4(!w15), .Z5(!Z5), .Z6(!w12), .Z7(!w10));   //: @(852,169) /sn:0 /w:[ 1 0 1 0 1 1 1 0 1 1 ]
  register R4 (.Q(w16), .D(DIN), .EN(w15), .CLR(w4), .CK(!w0));   //: @(531,358) /w:[ 0 27 0 13 21 ]
  //: joint g7 (R10) @(532, 600) /w:[ 2 -1 1 4 ]
  //: joint g22 (w4) @(586, 337) /w:[ 5 -1 6 12 ]
  //: joint g31 (w4) @(863, 417) /w:[ 17 -1 18 28 ]
  register R1 (.Q(R2), .D(DIN), .EN(w3), .CLR(w4), .CK(!w0));   //: @(262,449) /w:[ 5 21 1 23 11 ]
  register R3 (.Q(R3), .D(DIN), .EN(w7), .CLR(w4), .CK(!w0));   //: @(433,446) /w:[ 3 25 0 25 7 ]
  //: joint g33 (w4) @(673, 417) /w:[ 19 -1 20 26 ]
  //: joint g41 (DIN) @(717, 320) /w:[ 6 -1 5 8 ]
  //: joint g36 (w4) @(904, 337) /w:[ 1 -1 2 16 ]
  //: joint g40 (DIN) @(433, 320) /w:[ 13 -1 14 24 ]
  //: joint g42 (DIN) @(629, 320) /w:[ 4 -1 3 10 ]
  //: joint g12 (w0) @(479, 381) /w:[ 18 20 17 -1 ]
  //: input g28 (clr) @(1034,337) /sn:0 /R:2 /w:[ 1 ]
  //: input g34 (clk) @(53,398) /sn:0 /w:[ 1 ]
  mux g14 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SA), .Z(AOUT));   //: @(279,657) /sn:0 /w:[ 5 0 5 5 3 0 0 3 0 0 ] /ss:0 /do:0
  //: input g5 (RegWr) @(46,363) /sn:0 /w:[ 0 ]
  //: joint g11 (w0) @(293, 381) /w:[ 16 22 15 -1 ]
  //: joint g21 (w4) @(388, 337) /w:[ 7 -1 8 10 ]
  //: joint g19 (R0) @(255, 523) /w:[ 1 -1 2 4 ]
  //: input g20 (SD) @(780,138) /sn:0 /w:[ 0 ]
  //: joint g32 (w4) @(487, 417) /w:[ 21 -1 22 24 ]
  register R0 (.Q(R0), .D(DIN), .EN(w8), .CLR(w4), .CK(!w0));   //: @(181,362) /w:[ 3 19 0 9 25 ]
  //: input g0 (DIN) @(531,267) /sn:0 /R:3 /w:[ 0 ]
  //: joint g15 (R5) @(527, 586) /w:[ 2 -1 1 4 ]
  //: joint g38 (w0) @(577, 481) /w:[ 1 2 4 -1 ]
  //: joint g27 (w0) @(125, 381) /w:[ 14 24 26 13 ]
  mux g13 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SB), .Z(BOUT));   //: @(516,659) /sn:0 /w:[ 0 3 3 0 5 5 5 5 1 1 ] /ss:0 /do:0

endmodule

module main;    //: root_module
supply0 w16;    //: /sn:0 {0}(1775,47)(1775,61){1}
supply0 w37;    //: /sn:0 {0}(2209,82)(2209,105){1}
supply0 w14;    //: /sn:0 {0}(1571,430)(1571,409){1}
supply0 w11;    //: /sn:0 {0}(1479,218)(1460,218){1}
wire [31:0] w13;    //: /sn:0 {0}(1421,224)(1421,273){1}
//: {2}(1423,275)(1531,275)(1531,69)(1761,69){3}
//: {4}(1421,277)(1421,384)(1553,384){5}
wire [31:0] w34;    //: /sn:0 {0}(2915,371)(2855,371)(2855,520)(2601,520)(2601,327){1}
//: {2}(2603,325)(2711,325){3}
//: {4}(2599,325)(2507,325){5}
wire [31:0] w4;    //: /sn:0 {0}(2384,-7)(1839,-7)(1839,190)(1706,190){1}
//: {2}(1704,188)(1704,171){3}
//: {4}(1704,192)(1704,212){5}
//: {6}(1704,213)(1704,243){7}
//: {8}(1704,244)(1704,276){9}
//: {10}(1704,277)(1704,343){11}
//: {12}(1704,344)(1704,382)(1588,382){13}
wire w39;    //: /sn:0 {0}(2299,110)(2310,110)(2310,85){1}
wire w25;    //: /sn:0 {0}(1819,455)(2047,455)(2047,385){1}
wire w0;    //: /sn:0 {0}(1309,492)(1641,492){1}
//: {2}(1645,492)(1854,492)(1854,165)(1981,165)(1981,181){3}
//: {4}(1643,490)(1643,275){5}
wire [31:0] w22;    //: /sn:0 /dp:1 {0}(1610,129)(1610,139)(1724,139)(1724,101)(1761,101){1}
wire w20;    //: /sn:0 {0}(1985,418)(1996,418)(1996,385){1}
wire [31:0] w29;    //: /sn:0 {0}(2188,313)(2321,313){1}
wire [4:0] w30;    //: /sn:0 {0}(1864,277)(1708,277){1}
wire [31:0] w42;    //: /sn:0 {0}(2083,342)(2105,342){1}
//: {2}(2109,342)(2151,342)(2151,323)(2159,323){3}
//: {4}(2107,340)(2107,145)(2195,145){5}
wire w19;    //: /sn:0 {0}(1643,259)(1643,208)(1460,208){1}
wire [31:0] w18;    //: /sn:0 {0}(1790,85)(2150,85){1}
//: {2}(2152,83)(2152,52)(2294,52){3}
//: {4}(2152,87)(2152,113)(2195,113){5}
wire w23;    //: /sn:0 {0}(1793,312)(1864,312){1}
wire w21;    //: /sn:0 /dp:1 {0}(2209,172)(2209,153){1}
wire [3:0] w24;    //: /sn:0 /dp:1 {0}(2391,182)(2391,210){1}
wire w1;    //: /sn:0 {0}(1305,455)(1358,455){1}
//: {2}(1362,455)(1803,455){3}
//: {4}(1360,453)(1360,213)(1384,213){5}
wire [4:0] w31;    //: /sn:0 {0}(1864,244)(1708,244){1}
wire [4:0] w32;    //: /sn:0 /dp:1 {0}(1708,213)(1864,213){1}
wire w46;    //: /sn:0 {0}(2770,224)(2778,224)(2778,254){1}
wire w17;    //: /sn:0 {0}(2755,487)(2777,487)(2777,455){1}
wire [31:0] w44;    //: /sn:0 {0}(2323,62)(2344,62)(2344,13)(2384,13){1}
wire w33;    //: /sn:0 {0}(2909,407)(2931,407)(2931,384){1}
wire [31:0] w35;    //: /sn:0 /dp:1 {0}(2294,72)(2249,72)(2249,129)(2224,129){1}
wire [15:0] w28;    //: /sn:0 {0}(1864,344)(1708,344){1}
wire [31:0] w49;    //: /sn:0 {0}(2413,3)(2440,3)(2440,-52)(1421,-52)(1421,203){1}
wire [31:0] w45;    //: /sn:0 {0}(2083,213)(2214,213)(2214,249)(2321,249){1}
wire w2;    //: /sn:0 {0}(2169,369)(2175,369)(2175,336){1}
wire [31:0] w47;    //: /sn:0 {0}(2944,361)(2960,361)(2960,544)(1915,544)(1915,385){1}
wire w15;    //: /sn:0 /dp:1 {0}(2543,262)(2507,262){1}
wire w38;    //: /sn:0 {0}(2387,52)(2400,52)(2400,26){1}
wire [31:0] w43;    //: /sn:0 {0}(2836,351)(2915,351){1}
wire [31:0] w26;    //: /sn:0 {0}(2711,421)(2129,421)(2129,287){1}
//: {2}(2131,285)(2151,285)(2151,303)(2159,303){3}
//: {4}(2127,285)(2083,285){5}
wire w40;    //: /sn:0 /dp:1 {0}(1775,131)(1775,109){1}
//: enddecls

  //: switch g4 (w2) @(2152,369) /sn:0 /w:[ 0 ] /st:0
  MEM g44 (.MemWrite(w46), .Address(w34), .WriteData(w26), .MemRead(w17), .ReadData(w43));   //: @(2712, 255) /sz:(123, 199) /sn:0 /p:[ Ti0>1 Li0>3 Li1>0 Bi0>1 Ro0<0 ]
  //: joint g3 (w0) @(1643, 492) /w:[ 2 4 1 -1 ]
  //: switch g47 (w17) @(2738,487) /sn:0 /w:[ 0 ] /st:0
  register g16 (.Q(w13), .D(w49), .EN(w11), .CLR(w19), .CK(w1));   //: @(1421,213) /sn:0 /w:[ 0 1 1 1 5 ]
  //: switch g26 (w23) @(1776,312) /sn:0 /w:[ 0 ] /st:1
  //: supply0 g17 (w11) @(1485,218) /sn:0 /R:1 /w:[ 0 ]
  //: joint g2 (w1) @(1360, 455) /w:[ 2 4 1 -1 ]
  //: switch g30 (w20) @(1968,418) /sn:0 /w:[ 0 ] /st:1
  //: supply0 g23 (w16) @(1775,41) /sn:0 /R:2 /w:[ 0 ]
  clock g1 (.Z(w1));   //: @(1292,455) /sn:0 /w:[ 0 ] /omega:100 /phi:0 /duty:50
  mux g39 (.I0(w44), .I1(w4), .S(w38), .Z(w49));   //: @(2400,3) /sn:0 /R:1 /w:[ 1 0 1 0 ] /ss:0 /do:0
  READ g24 (.clr(w0), .Reg1(w32), .Reg2(w31), .RegMux(w30), .RegDst(w23), .ESignExt(w28), .Data(w47), .clk(w25), .RegWrite(w20), .Data1(w45), .SSignExt(w42), .Data2(w26));   //: @(1865, 182) /sz:(217, 202) /sn:0 /p:[ Ti0>3 Li0>1 Li1>0 Li2>0 Li3>1 Li4>0 Bi0>1 Bi1>1 Bi2>1 Ro0<0 Ro1<0 Ro2<5 ]
  tran g29(.Z(w31), .I(w4[20:16]));   //: @(1702,244) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  //: switch g51 (w38) @(2370,52) /sn:0 /w:[ 0 ] /st:0
  not g18 (.I(w0), .Z(w19));   //: @(1643,269) /sn:0 /R:1 /w:[ 5 0 ]
  tran g25(.Z(w32), .I(w4[25:21]));   //: @(1702,213) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  //: switch g49 (w33) @(2892,407) /sn:0 /w:[ 0 ] /st:0
  //: joint g50 (w34) @(2601, 325) /w:[ 2 -1 4 1 ]
  led g56 (.I(w21));   //: @(2209,179) /sn:0 /R:2 /w:[ 0 ] /type:0
  add g35 (.A(w42), .B(w18), .S(w35), .CI(w37), .CO(w21));   //: @(2211,129) /sn:0 /R:1 /w:[ 5 5 1 1 1 ]
  not g31 (.I(w1), .Z(w25));   //: @(1809,455) /sn:0 /w:[ 3 0 ]
  //: dip g22 (w22) @(1610,119) /sn:0 /w:[ 0 ] /st:1
  //: switch g45 (w46) @(2753,224) /sn:0 /w:[ 0 ] /st:0
  //: joint g41 (w4) @(1704, 190) /w:[ 1 2 -1 4 ]
  //: supply0 g36 (w37) @(2209,76) /sn:0 /R:2 /w:[ 0 ]
  ALU g33 (.ALUOp(w24), .B(w29), .A(w45), .Zero(w15), .ALURes(w34));   //: @(2322, 211) /sz:(184, 161) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Ro0<1 Ro1<5 ]
  //: switch g52 (w39) @(2282,110) /sn:0 /w:[ 0 ] /st:0
  //: joint g42 (w13) @(1421, 275) /w:[ 2 1 -1 4 ]
  //: joint g40 (w18) @(2152, 85) /w:[ -1 2 1 4 ]
  //: joint g46 (w26) @(2129, 285) /w:[ 2 -1 4 1 ]
  //: dip g34 (w24) @(2391,172) /sn:0 /w:[ 0 ] /st:0
  tran g28(.Z(w30), .I(w4[15:11]));   //: @(1702,277) /sn:0 /R:2 /w:[ 1 10 9 ] /ss:1
  rom g14 (.A(w13), .D(w4), .OE(w14));   //: @(1571,383) /sn:0 /w:[ 5 13 1 ]
  add g21 (.A(w22), .B(w13), .S(w18), .CI(w16), .CO(w40));   //: @(1777,85) /sn:0 /R:1 /w:[ 1 3 0 1 1 ]
  mux g32 (.I0(w42), .I1(w26), .S(w2), .Z(w29));   //: @(2175,313) /sn:0 /R:1 /w:[ 3 3 1 0 ] /ss:0 /do:0
  //: switch g0 (w0) @(1292,492) /sn:0 /w:[ 0 ] /st:0
  led g43 (.I(w15));   //: @(2550,262) /sn:0 /R:3 /w:[ 0 ] /type:0
  mux g38 (.I0(w18), .I1(w35), .S(w39), .Z(w44));   //: @(2310,62) /sn:0 /R:1 /w:[ 3 0 1 0 ] /ss:0 /do:1
  //: supply0 g15 (w14) @(1571,436) /sn:0 /w:[ 0 ]
  mux g48 (.I0(w34), .I1(w43), .S(w33), .Z(w47));   //: @(2931,361) /sn:0 /R:1 /w:[ 0 1 1 0 ] /ss:0 /do:0
  tran g27(.Z(w28), .I(w4[15:0]));   //: @(1702,344) /sn:0 /R:2 /w:[ 1 12 11 ] /ss:1
  //: joint g37 (w42) @(2107, 342) /w:[ 2 4 1 -1 ]
  led g55 (.I(w40));   //: @(1775,138) /sn:0 /R:2 /w:[ 0 ] /type:0

endmodule
