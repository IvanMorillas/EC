//: version "1.8.7"

module Sumador_HA(C, B, A, S);
//: interface  /sz:(183, 129) /bd:[ Li0>A(35/129) Li1>B(80/129) Ro0<S(62/129) Ro1<C(89/129) ]
input B;    //: /sn:0 {0}(354,174)(393,174)(393,173)(403,173){1}
//: {2}(407,173)(424,173)(424,159)(432,159){3}
//: {4}(405,175)(405,193)(429,193){5}
input A;    //: /sn:0 {0}(353,155)(380,155)(380,154)(390,154){1}
//: {2}(394,154)(432,154){3}
//: {4}(392,156)(392,188)(429,188){5}
output C;    //: /sn:0 {0}(515,191)(450,191){1}
output S;    //: /sn:0 {0}(515,157)(453,157){1}
//: enddecls

  //: output g4 (C) @(512,191) /sn:0 /w:[ 0 ]
  //: input g3 (B) @(352,174) /sn:0 /w:[ 0 ]
  //: input g2 (A) @(351,155) /sn:0 /w:[ 0 ]
  xor g1 (.I0(A), .I1(B), .Z(S));   //: @(443,157) /sn:0 /delay:" 4" /w:[ 3 3 1 ]
  //: joint g6 (A) @(392, 154) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(405, 173) /w:[ 2 -1 1 4 ]
  //: output g5 (S) @(512,157) /sn:0 /w:[ 0 ]
  and g0 (.I0(A), .I1(B), .Z(C));   //: @(440,191) /sn:0 /delay:" 3" /w:[ 5 5 1 ]

endmodule

module CPA(A, S, B, Cin);
//: interface  /sz:(114, 109) /bd:[ Ti0>A[3:0](80/114) Ti1>B[3:0](47/114) Ri0>Cin(36/109) Bo0<S[4:0](67/114) ]
input [3:0] B;    //: /sn:0 {0}(1157,146)(1089,146){1}
//: {2}(1088,146)(914,146){3}
//: {4}(913,146)(710,146){5}
//: {6}(709,146)(509,146){7}
//: {8}(508,146)(313,146){9}
input [3:0] A;    //: /sn:0 /dp:1 {0}(314,131)(469,131){1}
//: {2}(470,131)(696,131)(696,133){3}
//: {4}(696,134)(696,141)(879,141)(879,126)(894,126)(894,134){5}
//: {6}(894,135)(894,142)(965,142)(965,131)(1058,131){7}
//: {8}(1059,131)(1159,131){9}
input Cin;    //: /sn:0 {0}(1120,230)(1120,198)(1193,198){1}
output [4:0] S;    //: /sn:0 {0}(1397,420)(1250,420)(1250,425)(1240,425){1}
wire w6;    //: /sn:0 {0}(710,238)(710,150){1}
wire w13;    //: /sn:0 {0}(1106,339)(1106,360)(1006,360)(1006,213)(945,213)(945,231){1}
wire w16;    //: /sn:0 {0}(915,231)(915,158)(914,158)(914,150){1}
wire w7;    //: /sn:0 {0}(684,238)(684,134)(691,134){1}
wire w4;    //: /sn:0 {0}(479,329)(479,415)(1234,415){1}
wire w3;    //: /sn:0 {0}(526,329)(526,405)(1234,405){1}
wire w12;    //: /sn:0 {0}(1060,230)(1060,143)(1059,143)(1059,135){1}
wire w18;    //: /sn:0 {0}(930,333)(930,359)(838,359)(838,214)(756,214)(756,238){1}
wire w19;    //: /sn:0 {0}(887,333)(887,435)(1234,435){1}
wire w1;    //: /sn:0 {0}(509,237)(509,150){1}
wire w8;    //: /sn:0 {0}(739,330)(739,348)(625,348)(625,227)(543,227)(543,237){1}
wire w17;    //: /sn:0 {0}(881,231)(881,135)(889,135){1}
wire w14;    //: /sn:0 {0}(1066,339)(1066,445)(1234,445){1}
wire w2;    //: /sn:0 {0}(471,237)(471,143)(470,143)(470,135){1}
wire w11;    //: /sn:0 {0}(1091,230)(1091,158)(1089,158)(1089,150){1}
wire w9;    //: /sn:0 {0}(692,330)(692,425)(1234,425){1}
//: enddecls

  //: input g4 (A) @(312,131) /sn:0 /w:[ 0 ]
  tran g8(.Z(w2), .I(A[3]));   //: @(470,129) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: output g16 (S) @(1394,420) /sn:0 /w:[ 0 ]
  Sumador_FA g3 (.A(w17), .B(w16), .Cin(w13), .S(w19), .C(w18));   //: @(859, 232) /sz:(119, 100) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  Sumador_FA g2 (.A(w12), .B(w11), .Cin(Cin), .S(w14), .C(w13));   //: @(1040, 231) /sz:(110, 107) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Bo0<0 Bo1<0 ]
  Sumador_FA g1 (.A(w7), .B(w6), .Cin(w18), .S(w9), .C(w8));   //: @(660, 239) /sz:(132, 90) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  tran g10(.Z(w11), .I(B[0]));   //: @(1089,144) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g6(.Z(w17), .I(A[1]));   //: @(892,135) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:0
  tran g7(.Z(w7), .I(A[2]));   //: @(694,134) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:0
  //: input g9 (B) @(311,146) /sn:0 /w:[ 9 ]
  tran g12(.Z(w6), .I(B[2]));   //: @(710,144) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g5(.Z(w12), .I(A[0]));   //: @(1059,129) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g11(.Z(w16), .I(B[1]));   //: @(914,144) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: input g14 (Cin) @(1195,198) /sn:0 /R:2 /w:[ 1 ]
  concat g15 (.I0(w14), .I1(w19), .I2(w9), .I3(w4), .I4(w3), .Z(S));   //: @(1239,425) /sn:0 /w:[ 1 1 1 1 1 1 ] /dr:0
  Sumador_FA g0 (.A(w2), .B(w1), .Cin(w8), .S(w4), .C(w3));   //: @(447, 238) /sz:(133, 90) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  tran g13(.Z(w1), .I(B[3]));   //: @(509,144) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1

endmodule

module Sumador_FA(B, A, C, S, Cin);
//: interface  /sz:(90, 70) /bd:[ Li0>A(13/70) Li1>B(33/70) Li2>Cin(51/70) Ro0<S(17/70) Ro1<C(42/70) ]
input B;    //: /sn:0 {0}(67,222)(120,222)(120,219)(130,219){1}
input A;    //: /sn:0 /dp:1 {0}(69,193)(120,193)(120,194)(130,194){1}
input Cin;    //: /sn:0 {0}(71,286)(327,286)(327,261)(337,261){1}
output C;    //: /sn:0 {0}(574,310)(544,310)(544,309)(514,309){1}
output S;    //: /sn:0 /dp:1 {0}(443,251)(584,251)(584,253)(594,253){1}
wire w7;    //: /sn:0 {0}(443,266)(483,266)(483,306)(493,306){1}
wire w2;    //: /sn:0 {0}(213,209)(273,209)(273,236)(337,236){1}
wire w9;    //: /sn:0 /dp:1 {0}(493,311)(264,311)(264,224)(213,224){1}
//: enddecls

  //: input g4 (B) @(65,222) /sn:0 /w:[ 0 ]
  //: input g3 (A) @(67,193) /sn:0 /w:[ 0 ]
  or g2 (.I0(w7), .I1(w9), .Z(C));   //: @(504,309) /sn:0 /delay:" 3" /w:[ 1 0 1 ]
  Sumador_HA g1 (.B(Cin), .A(w2), .C(w7), .S(S));   //: @(338, 218) /sz:(104, 70) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: output g6 (C) @(571,310) /sn:0 /w:[ 0 ]
  //: output g7 (S) @(591,253) /sn:0 /w:[ 1 ]
  //: input g5 (Cin) @(69,286) /sn:0 /w:[ 0 ]
  Sumador_HA g0 (.B(B), .A(A), .C(w9), .S(w2));   //: @(131, 176) /sz:(81, 70) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]

endmodule

module main;    //: root_module
wire [15:0] w4;    //: /sn:0 {0}(540,261)(540,298)(622,298){1}
wire [15:0] w0;    //: /sn:0 {0}(495,290)(495,346)(622,346){1}
wire [15:0] w3;    //: /sn:0 {0}(950,288)(950,296)(913,296){1}
wire w1;    //: /sn:0 {0}(531,384)(622,384){1}
wire w2;    //: /sn:0 {0}(923,371)(913,371){1}
//: enddecls

  //: switch g3 (w1) @(514,384) /sn:0 /w:[ 0 ] /st:0
  //: dip g2 (w0) @(495,280) /sn:0 /w:[ 0 ] /st:0
  //: dip g1 (w4) @(540,251) /sn:0 /w:[ 0 ] /st:0
  CPA_Ex g0 (.Cin(w1), .B(w0), .A(w4), .Cout(w2), .S(w3));   //: @(623, 259) /sz:(289, 158) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Ro0<1 Ro1<1 ]

endmodule

module CPA_Ex(A, Cout, S, B, Cin);
//: interface  /sz:(289, 158) /bd:[ Li0>A[15:0](39/158) Li1>B[15:0](87/158) Li2>Cin(125/158) Ro0<S[15:0](37/158) Ro1<Cout(112/158) ]
input [15:0] B;    //: /sn:0 {0}(1189,92)(984,92){1}
//: {2}(983,92)(775,92){3}
//: {4}(774,92)(575,92){5}
//: {6}(574,92)(360,92){7}
//: {8}(359,92)(308,92){9}
input [15:0] A;    //: /sn:0 {0}(182,62)(392,62){1}
//: {2}(393,62)(577,62)(577,59){3}
//: {4}(577,58)(577,28)(824,28)(824,55){5}
//: {6}(824,56)(824,62)(1013,62){7}
//: {8}(1014,62)(1046,62){9}
input Cin;    //: /sn:0 {0}(1117,246)(1051,246){1}
output Cout;    //: /sn:0 /dp:1 {0}(375,352)(317,352)(317,448)(294,448){1}
output [15:0] S;    //: /sn:0 {0}(1312,449)(1139,449){1}
wire [3:0] w16;    //: /sn:0 {0}(803,454)(1133,454){1}
wire [3:0] w13;    //: /sn:0 {0}(360,96)(360,217){1}
wire w6;    //: /sn:0 {0}(998,341)(909,341)(909,251)(847,251){1}
wire [4:0] w7;    //: /sn:0 {0}(1003,471)(1003,465){1}
//: {2}(1003,464)(1003,341){3}
//: {4}(1003,340)(1003,320){5}
wire [3:0] w4;    //: /sn:0 {0}(819,56)(812,56)(812,214){1}
wire [3:0] w0;    //: /sn:0 {0}(1014,66)(1014,74)(1016,74)(1016,209){1}
wire [4:0] w20;    //: /sn:0 {0}(380,439)(380,433){1}
//: {2}(380,432)(380,352){3}
//: {4}(380,351)(380,328){5}
wire [3:0] w19;    //: /sn:0 {0}(1133,434)(389,434)(389,433)(384,433){1}
wire [3:0] w18;    //: /sn:0 {0}(1133,444)(599,444){1}
wire [3:0] w12;    //: /sn:0 {0}(393,66)(393,217){1}
wire w10;    //: /sn:0 {0}(794,360)(696,360)(696,251)(643,251){1}
wire [3:0] w1;    //: /sn:0 {0}(984,96)(984,104)(983,104)(983,209){1}
wire [3:0] w8;    //: /sn:0 {0}(581,59)(608,59)(608,214){1}
wire w14;    //: /sn:0 {0}(590,352)(497,352)(497,254)(428,254){1}
wire [3:0] w2;    //: /sn:0 /dp:1 {0}(1007,465)(1015,465)(1015,464)(1133,464){1}
wire [4:0] w11;    //: /sn:0 {0}(595,325)(595,351){1}
//: {2}(595,352)(595,443){3}
//: {4}(595,444)(595,449){5}
wire [4:0] w15;    //: /sn:0 {0}(799,459)(799,454){1}
//: {2}(799,453)(799,360){3}
//: {4}(799,359)(799,325){5}
wire [3:0] w5;    //: /sn:0 {0}(775,96)(775,104)(779,104)(779,214){1}
wire [3:0] w9;    //: /sn:0 {0}(575,96)(575,214){1}
//: enddecls

  tran g8(.Z(w12), .I(A[15:12]));   //: @(393,60) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: input g4 (A) @(180,62) /sn:0 /w:[ 0 ]
  tran g16(.Z(w10), .I(w15[4]));   //: @(797,360) /sn:0 /R:2 /anc:1 /w:[ 0 3 4 ] /ss:0
  CPA g3 (.B(w13), .A(w12), .Cin(w14), .S(w20));   //: @(313, 218) /sz:(114, 109) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<5 ]
  tran g17(.Z(w14), .I(w11[4]));   //: @(593,352) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:0
  CPA g2 (.B(w9), .A(w8), .Cin(w10), .S(w11));   //: @(528, 215) /sz:(114, 109) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<0 ]
  tran g23(.Z(w18), .I(w11[3:0]));   //: @(593,444) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  tran g24(.Z(w19), .I(w20[3:0]));   //: @(378,433) /sn:0 /R:2 /w:[ 1 1 2 ] /ss:1
  CPA g1 (.B(w5), .A(w4), .Cin(w6), .S(w15));   //: @(732, 215) /sz:(114, 109) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<5 ]
  //: output g18 (Cout) @(297,448) /sn:0 /R:2 /w:[ 1 ]
  //: output g25 (S) @(1309,449) /sn:0 /w:[ 0 ]
  tran g10(.Z(w1), .I(B[3:0]));   //: @(984,90) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  tran g6(.Z(w4), .I(A[7:4]));   //: @(822,56) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:0
  //: input g9 (B) @(1191,92) /sn:0 /R:2 /w:[ 0 ]
  tran g7(.Z(w8), .I(A[11:8]));   //: @(575,59) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:1
  tran g22(.Z(w16), .I(w15[3:0]));   //: @(797,454) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  tran g12(.Z(w9), .I(B[11:8]));   //: @(575,90) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  //: input g14 (Cin) @(1119,246) /sn:0 /R:2 /w:[ 0 ]
  tran g11(.Z(w5), .I(B[7:4]));   //: @(775,90) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  tran g5(.Z(w0), .I(A[3:0]));   //: @(1014,60) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g21(.Z(w2), .I(w7[3:0]));   //: @(1001,465) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  tran g19(.Z(Cout), .I(w20[4]));   //: @(378,352) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:0
  concat g20 (.I0(w2), .I1(w16), .I2(w18), .I3(w19), .Z(S));   //: @(1138,449) /sn:0 /w:[ 1 1 0 0 1 ] /dr:0
  tran g15(.Z(w6), .I(w7[4]));   //: @(1001,341) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:0
  CPA g0 (.B(w1), .A(w0), .Cin(Cin), .S(w7));   //: @(936, 210) /sz:(114, 109) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<5 ]
  tran g13(.Z(w13), .I(B[15:12]));   //: @(360,90) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1

endmodule
