//: version "1.8.7"

module CLL(G1, P3, P1, P0, G0, C2, P2, G3, C1, C4, G2, C3, C0);
//: interface  /sz:(818, 145) /bd:[ Ti0>G3(60/818) Ti1>P3(106/818) Ti2>G2(277/818) Ti3>P2(321/818) Ti4>P1(535/818) Ti5>G1(489/818) Ti6>P0(762/818) Ti7>G0(712/818) Ri0>C0(79/145) To0<C3(208/818) To1<C2(426/818) To2<C1(641/818) Lo0<C4(73/145) ]
input G2;    //: /sn:0 {0}(358,135)(358,326)(363,326){1}
//: {2}(367,326)(417,326)(417,330)(694,330){3}
//: {4}(365,328)(365,374)(384,374){5}
input C0;    //: /sn:0 {0}(466,132)(466,188)(514,188){1}
input P1;    //: /sn:0 {0}(377,134)(377,216)(452,216){1}
//: {2}(456,216)(520,216){3}
//: {4}(454,218)(454,226)(555,226){5}
output C3;    //: /sn:0 /dp:1 {0}(715,322)(769,322)(769,318)(821,318){1}
input G0;    //: /sn:0 /dp:5 {0}(445,132)(445,167){1}
//: {2}(447,169)(463,169)(463,178)(574,178){3}
//: {4}(445,171)(445,211)(520,211){5}
output C4;    //: /sn:0 /dp:1 {0}(774,376)(797,376)(797,374)(807,374){1}
output C2;    //: /sn:0 /dp:1 {0}(642,241)(736,241)(736,262)(815,262){1}
input P3;    //: /sn:0 /dp:11 {0}(505,373)(408,373)(408,363)(354,363)(354,369)(296,369){1}
//: {2}(294,367)(294,365)(293,365)(293,354){3}
//: {4}(295,352)(435,352)(435,362)(578,362){5}
//: {6}(293,350)(293,342){7}
//: {8}(295,340)(609,340)(609,357)(678,357){9}
//: {10}(293,338)(293,137){11}
//: {12}(294,371)(294,379)(384,379){13}
input G1;    //: /sn:0 {0}(401,133)(401,244){1}
//: {2}(403,246)(621,246){3}
//: {4}(401,248)(401,306)(446,306){5}
input G3;    //: /sn:0 {0}(317,137)(317,386)(753,386){1}
input P0;    //: /sn:0 {0}(425,130)(425,193)(514,193){1}
output C1;    //: /sn:0 /dp:1 {0}(595,181)(661,181)(661,218)(758,218)(758,245)(811,245){1}
input P2;    //: /sn:0 /dp:1 {0}(337,136)(337,264){1}
//: {2}(339,266)(572,266)(572,277)(602,277){3}
//: {4}(337,268)(337,276){5}
//: {6}(339,278)(466,278)(466,281)(523,281){7}
//: {8}(337,280)(337,311)(446,311){9}
wire w6;    //: /sn:0 {0}(576,229)(580,229){1}
//: {2}(584,229)(607,229)(607,241)(621,241){3}
//: {4}(582,231)(582,272)(602,272){5}
wire w7;    //: /sn:0 {0}(699,355)(745,355)(745,366)(753,366){1}
wire w3;    //: /sn:0 {0}(405,377)(455,377)(455,381)(753,381){1}
wire w18;    //: /sn:0 {0}(544,279)(571,279)(571,318){1}
//: {2}(573,320)(694,320){3}
//: {4}(569,320)(566,320)(566,357)(578,357){5}
wire w10;    //: /sn:0 {0}(526,371)(564,371)(564,376)(753,376){1}
wire w8;    //: /sn:0 {0}(623,275)(656,275)(656,278){1}
//: {2}(658,280)(686,280)(686,315)(694,315){3}
//: {4}(654,280)(649,280)(649,352)(678,352){5}
wire w2;    //: /sn:0 {0}(541,214)(543,214){1}
//: {2}(547,214)(614,214)(614,236)(621,236){3}
//: {4}(545,216)(545,261)(513,261)(513,276)(523,276){5}
wire w15;    //: /sn:0 {0}(467,309)(503,309)(503,323){1}
//: {2}(505,325)(694,325){3}
//: {4}(503,327)(503,368)(505,368){5}
wire w5;    //: /sn:0 {0}(535,191)(543,191)(543,190)(551,190){1}
//: {2}(555,190)(566,190)(566,183)(574,183){3}
//: {4}(553,192)(553,231)(555,231){5}
wire w9;    //: /sn:0 {0}(599,360)(647,360)(647,371)(753,371){1}
//: enddecls

  //: input g4 (G1) @(401,131) /sn:0 /R:3 /w:[ 0 ]
  //: input g8 (P3) @(293,135) /sn:0 /R:3 /w:[ 11 ]
  //: input g3 (P1) @(377,132) /sn:0 /R:3 /w:[ 0 ]
  and g16 (.I0(P1), .I1(w5), .Z(w6));   //: @(566,229) /sn:0 /w:[ 5 5 0 ]
  //: joint g26 (G1) @(401, 246) /w:[ 2 1 -1 4 ]
  //: joint g17 (G0) @(445, 169) /w:[ 2 1 -1 4 ]
  //: input g2 (P0) @(425,128) /sn:0 /R:3 /w:[ 0 ]
  //: joint g23 (w8) @(656, 280) /w:[ 2 1 4 -1 ]
  or g30 (.I0(w7), .I1(w9), .I2(w10), .I3(w3), .I4(G3), .Z(C4));   //: @(764,376) /sn:0 /w:[ 1 1 1 1 1 0 ]
  and g24 (.I0(G1), .I1(P2), .Z(w15));   //: @(457,309) /sn:0 /w:[ 5 9 0 ]
  and g39 (.I0(w8), .I1(P3), .Z(w7));   //: @(689,355) /sn:0 /w:[ 5 9 0 ]
  //: input g1 (G0) @(445,130) /sn:0 /R:3 /w:[ 0 ]
  //: joint g29 (P2) @(337, 278) /w:[ 6 5 -1 8 ]
  //: joint g18 (w5) @(553, 190) /w:[ 2 -1 1 4 ]
  and g25 (.I0(w2), .I1(P2), .Z(w18));   //: @(534,279) /sn:0 /w:[ 5 7 0 ]
  //: output g10 (C2) @(812,262) /sn:0 /w:[ 1 ]
  //: input g6 (P2) @(337,134) /sn:0 /R:3 /w:[ 0 ]
  //: joint g35 (P3) @(294, 369) /w:[ 1 2 -1 12 ]
  //: input g7 (G3) @(317,135) /sn:0 /R:3 /w:[ 0 ]
  //: output g9 (C1) @(808,245) /sn:0 /w:[ 1 ]
  and g22 (.I0(w6), .I1(P2), .Z(w8));   //: @(613,275) /sn:0 /w:[ 5 3 0 ]
  and g31 (.I0(G2), .I1(P3), .Z(w3));   //: @(395,377) /sn:0 /w:[ 5 13 0 ]
  //: joint g41 (w6) @(582, 229) /w:[ 2 -1 1 4 ]
  and g36 (.I0(w18), .I1(P3), .Z(w9));   //: @(589,360) /sn:0 /w:[ 5 5 0 ]
  and g33 (.I0(w15), .I1(P3), .Z(w10));   //: @(516,371) /sn:0 /w:[ 5 0 0 ]
  //: joint g40 (P3) @(293, 340) /w:[ 8 10 -1 7 ]
  //: output g12 (C4) @(804,374) /sn:0 /w:[ 1 ]
  //: joint g34 (w18) @(571, 320) /w:[ 2 1 4 -1 ]
  //: joint g28 (w2) @(545, 214) /w:[ 2 -1 1 4 ]
  //: input g5 (G2) @(358,133) /sn:0 /R:3 /w:[ 0 ]
  //: output g11 (C3) @(818,318) /sn:0 /w:[ 1 ]
  and g14 (.I0(C0), .I1(P0), .Z(w5));   //: @(525,191) /sn:0 /w:[ 1 1 0 ]
  or g21 (.I0(w8), .I1(w18), .I2(w15), .I3(G2), .Z(C3));   //: @(705,322) /sn:0 /w:[ 3 3 3 3 0 ]
  //: joint g19 (P1) @(454, 216) /w:[ 2 -1 1 4 ]
  //: joint g32 (G2) @(365, 326) /w:[ 2 -1 1 4 ]
  or g20 (.I0(w2), .I1(w6), .I2(G1), .Z(C2));   //: @(632,241) /sn:0 /w:[ 3 3 3 0 ]
  //: joint g38 (P2) @(337, 266) /w:[ 2 1 -1 4 ]
  //: input g0 (C0) @(466,130) /sn:0 /R:3 /w:[ 0 ]
  and g15 (.I0(G0), .I1(P1), .Z(w2));   //: @(531,214) /sn:0 /w:[ 5 3 0 ]
  //: joint g27 (w15) @(503, 325) /w:[ 2 1 -1 4 ]
  //: joint g37 (P3) @(293, 352) /w:[ 4 6 -1 3 ]
  or g13 (.I0(G0), .I1(w5), .Z(C1));   //: @(585,181) /sn:0 /w:[ 3 3 0 ]

endmodule

module PFA(Pi, Cin, B, S, Gi, A);
//: interface  /sz:(181, 159) /bd:[ Ti0>Cin(44/181) Ti1>B(106/181) Ti2>A(134/181) Bo0<Gi(49/181) Bo1<Pi(98/181) Bo2<S(129/181) ]
input B;    //: /sn:0 {0}(524,190)(573,190){1}
//: {2}(577,190)(698,190)(698,182)(708,182){3}
//: {4}(575,192)(575,273){5}
//: {6}(577,275)(688,275)(688,260)(800,260){7}
//: {8}(575,277)(575,288)(798,288){9}
output Gi;    //: /sn:0 /dp:1 {0}(819,291)(933,291){1}
input A;    //: /sn:0 {0}(526,152)(593,152){1}
//: {2}(597,152)(698,152)(698,177)(708,177){3}
//: {4}(595,154)(595,247){5}
//: {6}(597,249)(790,249)(790,255)(800,255){7}
//: {8}(595,251)(595,293)(798,293){9}
input Cin;    //: /sn:0 {0}(529,233)(770,233)(770,208)(802,208){1}
output Pi;    //: /sn:0 {0}(930,258)(821,258){1}
output S;    //: /sn:0 /dp:1 {0}(823,206)(930,206){1}
wire w2;    //: /sn:0 {0}(729,180)(792,180)(792,203)(802,203){1}
//: enddecls

  xor g4 (.I0(w2), .I1(Cin), .Z(S));   //: @(813,206) /sn:0 /delay:" 4" /w:[ 1 1 0 ]
  //: output g8 (Pi) @(927,258) /sn:0 /w:[ 0 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(719,180) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: input g2 (Cin) @(527,233) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(522,190) /sn:0 /w:[ 0 ]
  //: joint g10 (A) @(595, 152) /w:[ 2 -1 1 4 ]
  or g6 (.I0(A), .I1(B), .Z(Pi));   //: @(811,258) /sn:0 /delay:" 3" /w:[ 7 7 1 ]
  //: output g7 (S) @(927,206) /sn:0 /w:[ 1 ]
  //: output g9 (Gi) @(930,291) /sn:0 /w:[ 1 ]
  //: joint g12 (A) @(595, 249) /w:[ 6 5 -1 8 ]
  and g5 (.I0(B), .I1(A), .Z(Gi));   //: @(809,291) /sn:0 /delay:" 3" /w:[ 9 9 0 ]
  //: joint g11 (B) @(575, 190) /w:[ 2 -1 1 4 ]
  //: input g0 (A) @(524,152) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(575, 275) /w:[ 6 5 -1 8 ]

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 {0}(984,254)(984,244)(917,244){1}
wire w0;    //: /sn:0 {0}(722,405)(722,420)(714,420){1}
wire [3:0] w1;    //: /sn:0 {0}(837,405)(837,471)(826,471){1}
wire [3:0] w2;    //: /sn:0 /dp:1 {0}(698,172)(724,172)(724,210){1}
wire [3:0] w5;    //: /sn:0 /dp:1 {0}(800,169)(827,169)(827,210){1}
//: enddecls

  //: dip g4 (w2) @(660,172) /sn:0 /R:1 /w:[ 0 ] /st:8
  led g3 (.I(w1));   //: @(819,471) /sn:0 /R:1 /w:[ 1 ] /type:3
  //: switch g2 (w4) @(984,268) /sn:0 /R:1 /w:[ 0 ] /st:0
  led g1 (.I(w0));   //: @(707,420) /sn:0 /R:1 /w:[ 1 ] /type:0
  //: dip g5 (w5) @(762,169) /sn:0 /R:1 /w:[ 0 ] /st:7
  CLA g0 (.B(w2), .A(w5), .Cin(w4), .S(w1), .Cout(w0));   //: @(648, 211) /sz:(268, 193) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<0 Bo1<0 ]

endmodule

module CLA(A, S, Cout, Cin, B);
//: interface  /sz:(268, 193) /bd:[ Ti0>A[3:0](179/268) Ti1>B[3:0](76/268) Ri0>Cin(33/193) Bo0<Cout(74/268) Bo1<S[3:0](189/268) ]
input [3:0] B;    //: /sn:0 {0}(-161,-173)(-109,-173){1}
//: {2}(-108,-173)(116,-173){3}
//: {4}(117,-173)(330,-173){5}
//: {6}(331,-173)(542,-173){7}
//: {8}(543,-173)(654,-173){9}
input [3:0] A;    //: /sn:0 {0}(-159,-203)(-82,-203){1}
//: {2}(-81,-203)(143,-203){3}
//: {4}(144,-203)(252,-203)(252,-202)(359,-202){5}
//: {6}(360,-202)(465,-202)(465,-203)(568,-203){7}
//: {8}(569,-203)(650,-203){9}
input Cin;    //: /sn:0 /dp:1 {0}(481,48)(481,27)(737,27){1}
//: {2}(741,27)(841,27){3}
//: {4}(739,29)(739,420)(600,420){5}
output Cout;    //: /sn:0 {0}(-263,414)(-220,414){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(644,292)(682,292){1}
wire w16;    //: /sn:0 {0}(105,212)(105,330)(102,330)(102,340){1}
wire w13;    //: /sn:0 {0}(117,51)(117,-169){1}
wire w7;    //: /sn:0 {0}(331,45)(331,-169){1}
wire w22;    //: /sn:0 {0}(-117,213)(-117,330)(-113,330)(-113,340){1}
wire w36;    //: /sn:0 /dp:1 {0}(269,45)(269,35)(422,35)(422,340){1}
wire w0;    //: /sn:0 /dp:1 {0}(207,340)(207,41)(55,41)(55,51){1}
wire w3;    //: /sn:0 {0}(486,209)(486,330)(493,330)(493,340){1}
wire w20;    //: /sn:0 {0}(-81,52)(-81,-199){1}
wire w19;    //: /sn:0 {0}(-109,52)(-109,-161)(-108,-161)(-108,-169){1}
wire w12;    //: /sn:0 /dp:1 {0}(-11,340)(-11,42)(-171,42)(-171,52){1}
wire w23;    //: /sn:0 {0}(-86,213)(-86,277)(638,277){1}
wire w10;    //: /sn:0 {0}(323,206)(323,329)(316,329)(316,340){1}
wire w21;    //: /sn:0 {0}(-166,213)(-166,330)(-159,330)(-159,340){1}
wire w1;    //: /sn:0 {0}(543,48)(543,-169){1}
wire w8;    //: /sn:0 /dp:1 {0}(359,45)(359,-196)(360,-196)(360,-198){1}
wire w17;    //: /sn:0 {0}(140,212)(140,287)(638,287){1}
wire w14;    //: /sn:0 {0}(145,51)(145,-191)(144,-191)(144,-199){1}
wire w11;    //: /sn:0 {0}(354,206)(354,297)(638,297){1}
wire w2;    //: /sn:0 {0}(571,48)(571,-191)(569,-191)(569,-199){1}
wire w15;    //: /sn:0 {0}(60,212)(60,330)(58,330)(58,340){1}
wire w5;    //: /sn:0 {0}(566,209)(566,307)(638,307){1}
wire w26;    //: /sn:0 /dp:1 {0}(543,340)(543,330)(535,330)(535,209){1}
wire w9;    //: /sn:0 {0}(274,206)(274,330)(270,330)(270,340){1}
//: enddecls

  //: input g8 (A) @(-161,-203) /sn:0 /w:[ 0 ]
  CLL g4 (.G3(w21), .P3(w22), .G2(w15), .P2(w16), .P1(w10), .G1(w9), .P0(w26), .G0(w3), .C0(Cin), .C3(w12), .C2(w0), .C1(w36), .C4(Cout));   //: @(-219, 341) /sz:(818, 145) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>0 Ti7>1 Ri0>5 To0<0 To1<0 To2<1 Lo0<1 ]
  tran g16(.Z(w19), .I(B[3]));   //: @(-108,-175) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  PFA g3 (.A(w20), .B(w19), .Cin(w12), .S(w23), .Pi(w22), .Gi(w21));   //: @(-215, 53) /sz:(181, 159) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 Bo2<0 ]
  tran g17(.Z(w7), .I(B[1]));   //: @(331,-175) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  PFA g2 (.A(w14), .B(w13), .Cin(w0), .S(w17), .Pi(w16), .Gi(w15));   //: @(11, 52) /sz:(181, 159) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 Bo2<0 ]
  PFA g1 (.A(w8), .B(w7), .Cin(w36), .S(w11), .Pi(w10), .Gi(w9));   //: @(226, 46) /sz:(180, 159) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Bo0<0 Bo1<0 Bo2<0 ]
  //: output g18 (S) @(679,292) /sn:0 /w:[ 1 ]
  tran g10(.Z(w14), .I(A[2]));   //: @(144,-205) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: joint g6 (Cin) @(739, 27) /w:[ 2 -1 1 4 ]
  tran g9(.Z(w2), .I(A[0]));   //: @(569,-205) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: output g7 (Cout) @(-260,414) /sn:0 /R:2 /w:[ 0 ]
  tran g12(.Z(w8), .I(A[1]));   //: @(360,-204) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g14(.Z(w1), .I(B[0]));   //: @(543,-175) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g11(.Z(w20), .I(A[3]));   //: @(-81,-205) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: input g5 (Cin) @(843,27) /sn:0 /R:2 /w:[ 3 ]
  concat g19 (.I0(w5), .I1(w11), .I2(w17), .I3(w23), .Z(S));   //: @(643,292) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  tran g15(.Z(w13), .I(B[2]));   //: @(117,-175) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  PFA g0 (.A(w2), .B(w1), .Cin(Cin), .S(w5), .Pi(w26), .Gi(w3));   //: @(437, 49) /sz:(181, 159) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Bo0<0 Bo1<1 Bo2<0 ]
  //: input g13 (B) @(-163,-173) /sn:0 /w:[ 0 ]

endmodule
