//: version "1.8.7"

module Sumador_HA(C, B, A, S);
//: interface  /sz:(183, 129) /bd:[ Li0>A(35/129) Li1>B(80/129) Li2>B(80/129) Li3>A(35/129) Ro0<S(62/129) Ro1<C(89/129) Ro2<C(89/129) Ro3<S(62/129) ]
input B;    //: /sn:0 {0}(354,174)(393,174)(393,173)(403,173){1}
//: {2}(407,173)(424,173)(424,159)(432,159){3}
//: {4}(405,175)(405,193)(429,193){5}
input A;    //: /sn:0 {0}(353,155)(380,155)(380,154)(390,154){1}
//: {2}(394,154)(432,154){3}
//: {4}(392,156)(392,188)(429,188){5}
output C;    //: /sn:0 {0}(515,191)(450,191){1}
output S;    //: /sn:0 {0}(515,157)(453,157){1}
//: enddecls

  //: output g4 (C) @(512,191) /sn:0 /w:[ 0 ]
  //: input g3 (B) @(352,174) /sn:0 /w:[ 0 ]
  //: input g2 (A) @(351,155) /sn:0 /w:[ 0 ]
  xor g1 (.I0(A), .I1(B), .Z(S));   //: @(443,157) /sn:0 /delay:" 4" /w:[ 3 3 1 ]
  //: joint g6 (A) @(392, 154) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(405, 173) /w:[ 2 -1 1 4 ]
  //: output g5 (S) @(512,157) /sn:0 /w:[ 0 ]
  and g0 (.I0(A), .I1(B), .Z(C));   //: @(440,191) /sn:0 /delay:" 3" /w:[ 5 5 1 ]

endmodule

module CSA(Cout, A, S, B, Cin);
//: interface  /sz:(249, 190) /bd:[ Li0>A[3:0](41/190) Li1>B[3:0](89/190) Li2>Cin(144/190) Ro0<S[3:0](61/190) Ro1<Cout(129/190) ]
input [3:0] B;    //: /sn:0 /dp:1 {0}(686,180)(686,108){1}
//: {2}(688,106)(831,106)(831,181){3}
//: {4}(684,106)(683,106)(683,94)(487,94){5}
input [3:0] A;    //: /sn:0 {0}(469,61)(724,61)(724,69){1}
//: {2}(726,71)(867,71)(867,181){3}
//: {4}(724,73)(724,180){5}
input Cin;    //: /sn:0 /dp:1 {0}(425,198)(425,187)(309,187)(309,433)(359,433){1}
//: {2}(361,431)(361,365)(377,365){3}
//: {4}(361,435)(361,436)(733,436){5}
output Cout;    //: /sn:0 /dp:1 {0}(412,221)(349,221)(349,258)(359,258){1}
output [3:0] S;    //: /sn:0 {0}(756,449)(756,537)(794,537){1}
wire w4;    //: /sn:0 {0}(784,156)(799,156)(799,181){1}
wire [3:0] w3;    //: /sn:0 {0}(836,284)(836,401)(766,401)(766,420){1}
wire w0;    //: /sn:0 {0}(762,232)(504,232)(504,231)(441,231){1}
wire w18;    //: /sn:0 {0}(768,156)(758,156)(758,137)(664,137){1}
//: {2}(660,137)(482,137){3}
//: {4}(662,139)(662,149)(664,149)(664,180){5}
wire w2;    //: /sn:0 {0}(627,223)(606,223)(606,211)(441,211){1}
wire [3:0] w5;    //: /sn:0 /dp:1 {0}(746,420)(746,409)(680,409)(680,278){1}
//: enddecls

  //: output g8 (Cout) @(356,258) /sn:0 /w:[ 1 ]
  //: input g4 (A) @(467,61) /sn:0 /w:[ 0 ]
  mux g3 (.I0(w2), .I1(w0), .S(Cin), .Z(Cout));   //: @(425,221) /sn:0 /R:3 /delay:" 2 2" /w:[ 1 1 0 0 ] /ss:0 /do:0
  //: switch g16 (w18) @(465,137) /sn:0 /w:[ 3 ] /st:0
  //: joint g2 (w18) @(662, 137) /w:[ 1 -1 2 4 ]
  CPA g1 (.Cin(w4), .B(B), .A(A), .Cout(w0), .S(w3));   //: @(763, 182) /sz:(135, 101) /sn:0 /p:[ Ti0>1 Ti1>3 Ti2>3 Lo0<0 Bo0<0 ]
  //: output g10 (S) @(791,537) /sn:0 /w:[ 1 ]
  //: joint g6 (A) @(724, 71) /w:[ 2 1 -1 4 ]
  //: joint g7 (B) @(686, 106) /w:[ 2 -1 4 1 ]
  not g9 (.I(w18), .Z(w4));   //: @(774,156) /sn:0 /w:[ 0 0 ]
  mux g12 (.I0(w5), .I1(w3), .S(Cin), .Z(S));   //: @(756,436) /sn:0 /delay:" 2 2" /w:[ 0 1 5 0 ] /ss:0 /do:0
  //: input g11 (B) @(485,94) /sn:0 /w:[ 5 ]
  //: input g5 (Cin) @(379,365) /sn:0 /R:2 /w:[ 3 ]
  CPA g0 (.Cin(w18), .B(B), .A(A), .Cout(w2), .S(w5));   //: @(628, 181) /sz:(107, 96) /sn:0 /p:[ Ti0>5 Ti1>0 Ti2>5 Lo0<0 Bo0<1 ]
  //: joint g13 (Cin) @(361, 433) /w:[ -1 2 1 4 ]

endmodule

module CSA_16(S, Cin, B, Cout, A);
//: interface  /sz:(289, 164) /bd:[ Ti0>A[15:0](84/289) Ti1>B[15:0](170/289) Ti2>Cin(245/289) Bo0<S[15:0](98/289) Bo1<Cout(231/289) ]
input [15:0] B;    //: /sn:0 {0}(117,209)(205,209){1}
//: {2}(206,209)(352,209){3}
//: {4}(353,209)(486,209)(486,203){5}
//: {6}(486,202)(486,197)(596,197)(596,209)(717,209){7}
//: {8}(718,209)(725,209){9}
input [15:0] A;    //: /sn:0 {0}(117,179)(174,179){1}
//: {2}(175,179)(320,179){3}
//: {4}(321,179)(440,179)(440,174){5}
//: {6}(440,173)(440,169)(575,169)(575,179)(738,179){7}
//: {8}(739,179)(747,179){9}
input Cin;    //: /sn:0 /dp:1 {0}(759,350)(835,350){1}
output Cout;    //: /sn:0 {0}(249,428)(234,428)(234,418){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(846,526)(900,526)(900,532)(968,532){1}
wire [3:0] w6;    //: /sn:0 {0}(465,296)(465,174)(444,174){1}
wire w16;    //: /sn:0 {0}(840,491)(360,491)(360,477)(340,477){1}
wire w13;    //: /sn:0 {0}(840,521)(426,521)(426,525)(312,525){1}
wire w7;    //: /sn:0 {0}(840,581)(740,581){1}
wire w34;    //: /sn:0 {0}(381,419)(381,430)(288,430)(288,285)(245,285)(245,295){1}
wire [3:0] w25;    //: /sn:0 {0}(175,295)(175,183){1}
wire w4;    //: /sn:0 {0}(740,601)(840,601){1}
wire [3:0] w22;    //: /sn:0 {0}(758,620)(751,620){1}
//: {2}(750,620)(736,620)(736,601){3}
//: {4}(736,600)(736,592)(736,592)(736,581){5}
//: {6}(736,580)(736,569){7}
//: {8}(736,568)(736,399){9}
wire w3;    //: /sn:0 /dp:1 {0}(696,399)(696,409)(619,409)(619,286)(535,286)(535,296){1}
wire [3:0] w0;    //: /sn:0 {0}(739,183)(739,191)(740,191)(740,320){1}
wire w20;    //: /sn:0 {0}(193,445)(516,445)(516,451)(840,451){1}
wire [3:0] w30;    //: /sn:0 {0}(322,293)(322,191)(321,191)(321,183){1}
wire w19;    //: /sn:0 {0}(840,461)(175,461)(175,457){1}
wire w18;    //: /sn:0 {0}(840,471)(204,471)(204,469)(193,469){1}
wire w12;    //: /sn:0 {0}(840,531)(484,531)(484,523)(473,523){1}
wire [3:0] w23;    //: /sn:0 {0}(478,422)(478,511)(469,511)(469,522){1}
//: {2}(469,523)(469,533)(472,533)(472,540){3}
//: {4}(472,541)(472,547)(456,547)(456,564)(465,564){5}
//: {6}(466,564)(474,564)(474,584){7}
//: {8}(474,585)(474,590){9}
wire w10;    //: /sn:0 {0}(840,551)(466,551)(466,559){1}
wire w24;    //: /sn:0 {0}(525,422)(525,433)(430,433)(430,283)(392,283)(392,293){1}
wire [3:0] w21;    //: /sn:0 {0}(497,296)(497,203)(490,203){1}
wire [3:0] w31;    //: /sn:0 {0}(354,293)(354,221)(353,221)(353,213){1}
wire [3:0] w1;    //: /sn:0 {0}(718,213)(718,320){1}
wire w8;    //: /sn:0 {0}(840,571)(748,571)(748,569)(740,569){1}
wire w17;    //: /sn:0 {0}(840,481)(193,481){1}
wire [3:0] w33;    //: /sn:0 {0}(336,419)(336,476){1}
//: {2}(336,477)(336,492)(319,492){3}
//: {4}(318,492)(288,492)(288,506)(293,506){5}
//: {6}(294,506)(308,506)(308,524){7}
//: {8}(308,525)(308,531){9}
wire [3:0] w28;    //: /sn:0 /dp:3 {0}(189,418)(189,444){1}
//: {2}(189,445)(189,453)(175,453){3}
//: {4}(174,453)(156,453)(156,462)(189,462)(189,468){5}
//: {6}(189,469)(189,480){7}
//: {8}(189,481)(189,504){9}
wire w14;    //: /sn:0 {0}(840,511)(319,511)(319,496){1}
wire w11;    //: /sn:0 {0}(840,541)(476,541){1}
wire w15;    //: /sn:0 /dp:1 {0}(840,501)(294,501)(294,501){1}
wire w5;    //: /sn:0 {0}(751,615)(751,591)(840,591){1}
wire [3:0] w26;    //: /sn:0 {0}(207,295)(207,221)(206,221)(206,213){1}
wire w9;    //: /sn:0 {0}(840,561)(486,561)(486,585)(478,585){1}
//: enddecls

  tran g8(.Z(w5), .I(w22[1]));   //: @(751,618) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:0
  //: output g4 (S) @(965,532) /sn:0 /w:[ 1 ]
  tran g16(.Z(w12), .I(w23[3]));   //: @(467,523) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  //: input g3 (Cin) @(837,350) /sn:0 /R:2 /w:[ 1 ]
  tran g26(.Z(w0), .I(A[3:0]));   //: @(739,177) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g17(.Z(w13), .I(w33[0]));   //: @(306,525) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  CPA g2 (.B(w1), .A(w0), .Cin(Cin), .Cout(w3), .S(w22));   //: @(672, 321) /sz:(86, 77) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<9 ]
  tran g30(.Z(w31), .I(B[11:8]));   //: @(353,207) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g23(.Z(w19), .I(w28[2]));   //: @(175,451) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g24(.Z(w20), .I(w28[3]));   //: @(187,445) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: input g1 (B) @(115,209) /sn:0 /w:[ 0 ]
  tran g29(.Z(w21), .I(B[7:4]));   //: @(484,203) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:1
  tran g18(.Z(w14), .I(w33[1]));   //: @(319,490) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g25(.Z(w15), .I(w33[2]));   //: @(294,504) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:0
  CSA g10 (.Cin(w3), .B(w21), .A(w6), .Cout(w24), .S(w23));   //: @(437, 297) /sz:(130, 124) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<0 ]
  tran g6(.Z(w4), .I(w22[0]));   //: @(734,601) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:1
  tran g9(.Z(w8), .I(w22[3]));   //: @(734,569) /sn:0 /R:2 /w:[ 1 7 8 ] /ss:1
  tran g7(.Z(w7), .I(w22[2]));   //: @(734,581) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:1
  tran g31(.Z(w30), .I(A[11:8]));   //: @(321,177) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g22(.Z(w18), .I(w28[1]));   //: @(187,469) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  tran g33(.Z(w25), .I(A[15:12]));   //: @(175,177) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  CSA g12 (.Cin(w24), .B(w31), .A(w30), .Cout(w34), .S(w33));   //: @(295, 294) /sz:(128, 124) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<0 ]
  tran g28(.Z(w6), .I(A[7:4]));   //: @(438,174) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:1
  tran g14(.Z(w11), .I(w23[2]));   //: @(470,541) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  CSA g11 (.Cin(w34), .B(w26), .A(w25), .Cout(Cout), .S(w28));   //: @(148, 296) /sz:(128, 121) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<1 Bo1<0 ]
  concat g5 (.I0(w4), .I1(w5), .I2(w7), .I3(w8), .I4(w9), .I5(w10), .I6(w11), .I7(w12), .I8(w13), .I9(w14), .I10(w15), .I11(w16), .I12(w17), .I13(w18), .I14(w19), .I15(w20), .Z(S));   //: @(845,526) /sn:0 /w:[ 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 ] /dr:0
  tran g21(.Z(w17), .I(w28[0]));   //: @(187,481) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  tran g19(.Z(w16), .I(w33[3]));   //: @(334,477) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  tran g32(.Z(w26), .I(B[15:12]));   //: @(206,207) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: output g20 (Cout) @(246,428) /sn:0 /w:[ 0 ]
  tran g15(.Z(w10), .I(w23[1]));   //: @(466,562) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:0
  //: input g0 (A) @(115,179) /sn:0 /w:[ 0 ]
  tran g27(.Z(w1), .I(B[3:0]));   //: @(718,207) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g13(.Z(w9), .I(w23[0]));   //: @(472,585) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1

endmodule

module CPA(A, S, Cout, B, Cin);
//: interface  /sz:(86, 77) /bd:[ Ti0>A[3:0](68/86) Ti1>B[3:0](46/86) Ri0>Cin(29/77) Bo0<S[3:0](64/86) Bo1<Cout(24/86) ]
input [3:0] B;    //: /sn:0 {0}(1157,146)(1089,146){1}
//: {2}(1088,146)(914,146){3}
//: {4}(913,146)(710,146){5}
//: {6}(709,146)(509,146){7}
//: {8}(508,146)(313,146){9}
input [3:0] A;    //: /sn:0 /dp:1 {0}(314,131)(469,131){1}
//: {2}(470,131)(696,131)(696,133){3}
//: {4}(696,134)(696,141)(879,141)(879,126)(894,126)(894,134){5}
//: {6}(894,135)(894,142)(965,142)(965,131)(1058,131){7}
//: {8}(1059,131)(1159,131){9}
input Cin;    //: /sn:0 {0}(1120,230)(1120,198)(1193,198){1}
output Cout;    //: /sn:0 /dp:1 {0}(526,329)(526,458)(560,458){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(1397,420)(1250,420)(1250,425)(1240,425){1}
wire w16;    //: /sn:0 {0}(915,231)(915,158)(914,158)(914,150){1}
wire w13;    //: /sn:0 {0}(1106,339)(1106,360)(1006,360)(1006,213)(945,213)(945,231){1}
wire w6;    //: /sn:0 {0}(710,238)(710,150){1}
wire w7;    //: /sn:0 {0}(684,238)(684,134)(691,134){1}
wire w4;    //: /sn:0 {0}(479,329)(479,410)(1234,410){1}
wire w19;    //: /sn:0 {0}(887,333)(887,430)(1234,430){1}
wire w18;    //: /sn:0 {0}(930,333)(930,359)(838,359)(838,214)(756,214)(756,238){1}
wire w12;    //: /sn:0 {0}(1060,230)(1060,143)(1059,143)(1059,135){1}
wire w1;    //: /sn:0 {0}(509,237)(509,150){1}
wire w8;    //: /sn:0 {0}(739,330)(739,348)(625,348)(625,227)(543,227)(543,237){1}
wire w17;    //: /sn:0 {0}(881,231)(881,135)(889,135){1}
wire w14;    //: /sn:0 {0}(1066,339)(1066,440)(1234,440){1}
wire w11;    //: /sn:0 {0}(1091,230)(1091,158)(1089,158)(1089,150){1}
wire w2;    //: /sn:0 {0}(471,237)(471,143)(470,143)(470,135){1}
wire w9;    //: /sn:0 {0}(692,330)(692,420)(1234,420){1}
//: enddecls

  tran g8(.Z(w2), .I(A[3]));   //: @(470,129) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: input g4 (A) @(312,131) /sn:0 /w:[ 0 ]
  Sumador_FA g3 (.A(w17), .B(w16), .Cin(w13), .S(w19), .C(w18));   //: @(859, 232) /sz:(119, 100) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  //: output g16 (S) @(1394,420) /sn:0 /w:[ 0 ]
  //: output g17 (Cout) @(557,458) /sn:0 /w:[ 1 ]
  Sumador_FA g2 (.A(w12), .B(w11), .Cin(Cin), .S(w14), .C(w13));   //: @(1040, 231) /sz:(110, 107) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Bo0<0 Bo1<0 ]
  Sumador_FA g1 (.A(w7), .B(w6), .Cin(w18), .S(w9), .C(w8));   //: @(660, 239) /sz:(132, 90) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  tran g10(.Z(w11), .I(B[0]));   //: @(1089,144) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g6(.Z(w17), .I(A[1]));   //: @(892,135) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:0
  //: input g9 (B) @(311,146) /sn:0 /w:[ 9 ]
  tran g7(.Z(w7), .I(A[2]));   //: @(694,134) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:0
  tran g12(.Z(w6), .I(B[2]));   //: @(710,144) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: input g14 (Cin) @(1195,198) /sn:0 /R:2 /w:[ 1 ]
  tran g11(.Z(w16), .I(B[1]));   //: @(914,144) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g5(.Z(w12), .I(A[0]));   //: @(1059,129) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  Sumador_FA g0 (.A(w2), .B(w1), .Cin(w8), .S(w4), .C(Cout));   //: @(447, 238) /sz:(133, 90) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  concat g15 (.I0(w14), .I1(w19), .I2(w9), .I3(w4), .Z(S));   //: @(1239,425) /sn:0 /w:[ 1 1 1 1 1 ] /dr:0
  tran g13(.Z(w1), .I(B[3]));   //: @(509,144) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1

endmodule

module Sumador_FA(B, A, C, S, Cin);
//: interface  /sz:(90, 70) /bd:[ Li0>A(13/70) Li1>B(33/70) Li2>Cin(51/70) Li3>Cin(51/70) Li4>B(33/70) Li5>A(13/70) Ro0<S(17/70) Ro1<C(42/70) Ro2<C(42/70) Ro3<S(17/70) ]
input B;    //: /sn:0 {0}(67,222)(120,222)(120,219)(130,219){1}
input A;    //: /sn:0 /dp:1 {0}(69,193)(120,193)(120,194)(130,194){1}
input Cin;    //: /sn:0 {0}(71,286)(327,286)(327,261)(337,261){1}
output C;    //: /sn:0 {0}(574,310)(544,310)(544,309)(514,309){1}
output S;    //: /sn:0 /dp:1 {0}(443,251)(584,251)(584,253)(594,253){1}
wire w7;    //: /sn:0 {0}(443,266)(483,266)(483,306)(493,306){1}
wire w2;    //: /sn:0 {0}(213,209)(273,209)(273,236)(337,236){1}
wire w9;    //: /sn:0 /dp:1 {0}(493,311)(264,311)(264,224)(213,224){1}
//: enddecls

  //: input g4 (B) @(65,222) /sn:0 /w:[ 0 ]
  //: input g3 (A) @(67,193) /sn:0 /w:[ 0 ]
  or g2 (.I0(w7), .I1(w9), .Z(C));   //: @(504,309) /sn:0 /delay:" 3" /w:[ 1 0 1 ]
  Sumador_HA g1 (.B(Cin), .A(w2), .C(w7), .S(S));   //: @(338, 218) /sz:(104, 70) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: output g6 (C) @(571,310) /sn:0 /w:[ 0 ]
  //: output g7 (S) @(591,253) /sn:0 /w:[ 1 ]
  //: input g5 (Cin) @(69,286) /sn:0 /w:[ 0 ]
  Sumador_HA g0 (.B(B), .A(A), .C(w9), .S(w2));   //: @(131, 176) /sz:(81, 70) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 {0}(689,403)(689,443)(701,443){1}
wire [15:0] w3;    //: /sn:0 {0}(556,403)(556,524)(477,524)(477,503){1}
wire [15:0] w0;    //: /sn:0 {0}(484,129)(484,201)(542,201)(542,237){1}
wire [15:0] w1;    //: /sn:0 /dp:1 {0}(581,130)(581,221)(628,221)(628,237){1}
wire w2;    //: /sn:0 {0}(688,182)(703,182)(703,237){1}
//: enddecls

  led g4 (.I(w3));   //: @(477,496) /sn:0 /w:[ 1 ] /type:3
  //: switch g3 (w2) @(671,182) /sn:0 /w:[ 0 ] /st:0
  //: dip g2 (w1) @(581,120) /sn:0 /w:[ 0 ] /st:0
  //: dip g1 (w0) @(484,119) /sn:0 /w:[ 0 ] /st:0
  led g5 (.I(w4));   //: @(708,443) /sn:0 /R:3 /w:[ 1 ] /type:0
  CSA_16 g0 (.Cin(w2), .B(w1), .A(w0), .Cout(w4), .S(w3));   //: @(458, 238) /sz:(289, 164) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Bo0<0 Bo1<0 ]

endmodule
